
module ELM_inference_engine_tb;
    parameter input_cnt=10;//number of test inputs (which are stored in the X_test.txt file)
    reg clk,rst,start; // If rst = 1-->system will reset, if start=1 (rst=0): testing process starts,  
    reg din; //Test input
    reg din_valid; //If din_valid = 1 : Test Data which is to fed is still available ; else : Test_data = 0 : No test data to process (System remains idle) : state7    
    wire give_input; // Input is fed into the ELM inference engine if give_input=1 
    wire [3:0]hw_digit;//Decimal output
    wire output_valid; //Output is valid if output_valid = 1
    
    //Instantiating Inference engine
    ELM_inference_engine dm1(clk,rst,start,din,din_valid,give_input,hw_digit,output_valid);
  
     
    //initializing
    initial begin
        clk=0;rst=1;start=0;din_valid=1;
        #320 rst=0;start=1;
    end
    
    integer input_part,input_index,out_disp,display_done;
    reg [1:256]X_test[1:input_cnt];//Data memory (Test data : For test data storage [ Each row corresponds to a test vector (of 8 columns(each column=32bits)]-->256 bit input)  
    reg [3:0]Ytest_input[1:input_cnt];//Test outputs from "Y_test.txt" file : for comparison
    reg [3:0]Ytest_predict[1:input_cnt];//decimal outputs of all the test inputs
    reg [8:0]success;//9 bits for success (assuming max test inputs =493)

    initial begin
        input_part=1;input_index=1;success=0;display_done=0;//initialize the X_test array indices
        X_test[1] =256'b0000001111111100000001111000111000011110000001110011110000000111011110000000001111111000000000111111000000000011111100000000001111000000000000111100000000000111111000000000111011100000000011100110000000011100011110001111100000111111111000000001111110000000;
        X_test[2] =256'b0000000000000111000000000000111100000000001111000000000001111000000000011110000000000111111000000000111111000000001111111000000011111111000000000000111000000000000111000000000000111000000000000111000000000000011100000000000001100000000000000111000000000000;
        X_test[3] =256'b0111111100000000111000110000000011110011000000000011011100000000000001100000000000001110000000000000110000000000000110000000000000110000000000000111000000000000011000000000000001100000000000000110000000000000011000000000000001111111111111110001111111111000;
        X_test[4] =256'b1111111111111000000000000001100000000000000110000000000011110000000000111100000000000111100000000000111111111110000000000000001100000000000000110000000000000011000000000000011000000000000011100000000000111100000111000111000000011111111000000000111110000000;
        X_test[5] =256'b0000000000011111000000000011111000000000111110000000000111100000000000111000000000001111000000000001111000000000001110000000000001111000000000001110000000001100111111111111111011111111000011100000000000001110000000000000111000000000000011100000000000011110; 
        X_test[6] =256'b0000011111111100011111111000000011000000000000001100000000000000111000000000000001111000000000000001111100000000000000111111000000000000001111000000000000000111000000000000001100100000000000110111110000000011011111000000011100011111111111100000000001110000;
        X_test[7] =256'b0000000001111000000000001110000000000111110000000000111100000000000011100000000000111100000000000011100000000000011110000000000011111111111110001111000000111100111000000000111011100000000000111110000000000011111100000001111101111111111110000001111111100000;
        X_test[8] =256'b0000000000001111110000000011111001111111111110000011111101110000000000001110000000000000111000000000000111000000000000011000000000000011100000001111111111110000100001111111110000001110000011100000110000000000000011000000000000001100000000000000110000000000;
        X_test[9] =256'b0000011111111100000111110000111001111100000001110111100000000111001111000000111100011100000111100000111101111100000001111111000000111111110000000111111110000000111000011100000011000001111000001110000111100000011000011110000001111111110000000001111100000000;
        X_test[10]=256'b0011111110000000111110111111100011100000111111111100000000001111111000000011111111100000001111110111110000111111000111111111111000000111110011100000000000001110000000000000111100000000000001100000000000000111000000000000011100000000000001110000000000000111;
		  
        Ytest_input[1]=4'd0;Ytest_input[2]=4'd1;Ytest_input[3]=4'd2;Ytest_input[4]=4'd3;Ytest_input[5]=4'd4;
	Ytest_input[6]=4'd5;Ytest_input[7]=4'd6;Ytest_input[8]=4'd7;Ytest_input[9]=4'd8;Ytest_input[10]=4'd9;
    end
    always@(posedge clk)begin
        if(output_valid)begin //Indicates the Output of given test input vector is available
            if(hw_digit==Ytest_input[input_index])
                success=success+1;//success rate
            Ytest_predict[input_index]=hw_digit;//store decimal outputs
            input_index=input_index+1;input_part=1;//increasing the X_test array indices
        end

        if(input_index==input_cnt+1)begin //If all the test input vectors are given , then activate this signal : indicates there is No test input to process  
            din_valid=0;        
            if(display_done==0)begin
                $display("Given number and Predicted numbers :\n");
                for (out_disp=1;out_disp<=10;out_disp=out_disp+1)begin
                    $display("Input_digit = %d  , Predicted_digit = %d",Ytest_input[out_disp],Ytest_predict[out_disp]);
                end
                display_done=1;
           end
        end
        
        if(give_input)begin //pass the test input vector : if give_input=1 (Input is fed into design in 8 clock cycles)
            din=X_test[input_index][input_part];//send input part wise to design
            input_part=input_part+1;
        end
    end
    always #5 clk <= ~clk; 
endmodule