
module w21rom(clk,addr,d); 
    input clk;
    input [8:0] addr; // This is the 9 bit row address
    output reg [159:0] d; // data output of ROM : Entire row.

    wire [159:0] d_next ; // Declare as the wire. 
    wire [15:0]loc[1:420][1:10] ; // ROM organized as 256x420    
    reg [159:0]W21 ; // ROM organized as 256x420 

    //store Weights in temporary locations
    assign loc[1][1]=16'h0000,loc[1][2]=16'h0000,loc[1][3]=16'h0000,loc[1][4]=16'h0000,loc[1][5]=16'h0000,loc[1][6]=16'h0000,loc[1][7]=16'h0000,loc[1][8]=16'h0000,loc[1][9]=16'h0000,loc[1][10]=16'h0000,loc[2][1]=16'h0000,loc[2][2]=16'h0000,loc[2][3]=16'hffff,loc[2][4]=16'h0009,loc[2][5]=16'h0000,loc[2][6]=16'hfffd,loc[2][7]=16'h0006,loc[2][8]=16'hfffb,loc[2][9]=16'hfff4,loc[2][10]=16'h0005,loc[3][1]=16'hfffc,loc[3][2]=16'hffff,loc[3][3]=16'h0008,loc[3][4]=16'h0006,loc[3][5]=16'h000b,loc[3][6]=16'hffff,loc[3][7]=16'hfff8,loc[3][8]=16'hfff9,loc[3][9]=16'h0007,loc[3][10]=16'hfff5,loc[4][1]=16'h0005,loc[4][2]=16'h000a,loc[4][3]=16'hfffb,loc[4][4]=16'h0002,loc[4][5]=16'h0000,loc[4][6]=16'hfff7,loc[4][7]=16'h0002,loc[4][8]=16'hfff9,loc[4][9]=16'h0008,loc[4][10]=16'hfff5,loc[5][1]=16'hfffa,loc[5][2]=16'hffff,loc[5][3]=16'hfff6,loc[5][4]=16'h0002,loc[5][5]=16'hfffb,loc[5][6]=16'h0000,loc[5][7]=16'h0006,loc[5][8]=16'h0008,loc[5][9]=16'h0008,loc[5][10]=16'hfffb,loc[6][1]=16'hfffb,loc[6][2]=16'hfffb,loc[6][3]=16'h0001,loc[6][4]=16'h0001,loc[6][5]=16'h0000,loc[6][6]=16'h0005,loc[6][7]=16'hffff,loc[6][8]=16'h0002,loc[6][9]=16'hffff,loc[6][10]=16'h0004,loc[7][1]=16'h0002,loc[7][2]=16'h0005,loc[7][3]=16'h0001,loc[7][4]=16'h0002,loc[7][5]=16'h0001,loc[7][6]=16'h0001,loc[7][7]=16'h0000,loc[7][8]=16'h0000,loc[7][9]=16'h0004,loc[7][10]=16'hfff2,loc[8][1]=16'h000b,loc[8][2]=16'hffef,loc[8][3]=16'h0000,loc[8][4]=16'h0008,loc[8][5]=16'hfffa,loc[8][6]=16'hfffb,loc[8][7]=16'h0003,loc[8][8]=16'h000a,loc[8][9]=16'hfff7,loc[8][10]=16'h0007,loc[9][1]=16'h0007,loc[9][2]=16'hfff7,loc[9][3]=16'hfffb,loc[9][4]=16'h0003,loc[9][5]=16'h000a,loc[9][6]=16'hfff8,loc[9][7]=16'h0002,loc[9][8]=16'h0010,loc[9][9]=16'hfffe,loc[9][10]=16'hfff9,loc[10][1]=16'h0000,loc[10][2]=16'hfffb,loc[10][3]=16'h0002,loc[10][4]=16'h0005,loc[10][5]=16'h0000,loc[10][6]=16'h0000,loc[10][7]=16'hffff,loc[10][8]=16'h0008,loc[10][9]=16'hfff8,loc[10][10]=16'h0003,loc[11][1]=16'h0000,loc[11][2]=16'hfffc,loc[11][3]=16'hfffb,loc[11][4]=16'h0008,loc[11][5]=16'hfffc,loc[11][6]=16'hffff,loc[11][7]=16'h0001,loc[11][8]=16'hfffc,loc[11][9]=16'h0008,loc[11][10]=16'h0002,loc[12][1]=16'h0001,loc[12][2]=16'h0002,loc[12][3]=16'h0002,loc[12][4]=16'hfff1,loc[12][5]=16'h0003,loc[12][6]=16'h0008,loc[12][7]=16'hffff,loc[12][8]=16'h0005,loc[12][9]=16'h0000,loc[12][10]=16'hffff,loc[13][1]=16'h0001,loc[13][2]=16'h0003,loc[13][3]=16'h0006,loc[13][4]=16'hfffc,loc[13][5]=16'hfff7,loc[13][6]=16'h0000,loc[13][7]=16'hfffe,loc[13][8]=16'h0008,loc[13][9]=16'hfffe,loc[13][10]=16'h0001,loc[14][1]=16'hfffd,loc[14][2]=16'h000b,loc[14][3]=16'hfffc,loc[14][4]=16'h0007,loc[14][5]=16'hfffd,loc[14][6]=16'h0006,loc[14][7]=16'h0005,loc[14][8]=16'hffee,loc[14][9]=16'h0006,loc[14][10]=16'hfffa,loc[15][1]=16'hfffc,loc[15][2]=16'h0003,loc[15][3]=16'h0004,loc[15][4]=16'hfffa,loc[15][5]=16'h0001,loc[15][6]=16'hfffd,loc[15][7]=16'hfffb,loc[15][8]=16'h000c,loc[15][9]=16'hfffe,loc[15][10]=16'h0004,loc[16][1]=16'h0007,loc[16][2]=16'h0001,loc[16][3]=16'hfffe,loc[16][4]=16'h0001,loc[16][5]=16'h0000,loc[16][6]=16'h0001,loc[16][7]=16'hfffa,loc[16][8]=16'h0002,loc[16][9]=16'h0000,loc[16][10]=16'hfffd,loc[17][1]=16'hfffe,loc[17][2]=16'hfffd,loc[17][3]=16'h0006,loc[17][4]=16'h0001,loc[17][5]=16'h0005,loc[17][6]=16'hfff8,loc[17][7]=16'h000e,loc[17][8]=16'hfff7,loc[17][9]=16'hfff8,loc[17][10]=16'h0009,loc[18][1]=16'h0006,loc[18][2]=16'h0010,loc[18][3]=16'h0010,loc[18][4]=16'hfff3,loc[18][5]=16'h000d,loc[18][6]=16'h0002,loc[18][7]=16'hfff7,loc[18][8]=16'hffed,loc[18][9]=16'h0001,loc[18][10]=16'hfffb,loc[19][1]=16'h000a,loc[19][2]=16'hfffb,loc[19][3]=16'hfffe,loc[19][4]=16'h0002,loc[19][5]=16'hfffc,loc[19][6]=16'hfffc,loc[19][7]=16'hfff0,loc[19][8]=16'h0011,loc[19][9]=16'h000b,loc[19][10]=16'hfffd,loc[20][1]=16'hffff,loc[20][2]=16'h0003,loc[20][3]=16'hfff2,loc[20][4]=16'h0003,loc[20][5]=16'hfff9,loc[20][6]=16'h0004,loc[20][7]=16'h0010,loc[20][8]=16'h0009,loc[20][9]=16'h0003,loc[20][10]=16'hffee,loc[21][1]=16'h0001,loc[21][2]=16'h0003,loc[21][3]=16'h0003,loc[21][4]=16'hfffd,loc[21][5]=16'hfff9,loc[21][6]=16'h000a,loc[21][7]=16'h0001,loc[21][8]=16'h0009,loc[21][9]=16'hfff8,loc[21][10]=16'hfff9,loc[22][1]=16'hfff3,loc[22][2]=16'h0003,loc[22][3]=16'hfffe,loc[22][4]=16'hffff,loc[22][5]=16'h000e,loc[22][6]=16'h0007,loc[22][7]=16'hfffb,loc[22][8]=16'hfffd,loc[22][9]=16'h0008,loc[22][10]=16'hffff,loc[23][1]=16'h0000,loc[23][2]=16'h0000,loc[23][3]=16'h000a,loc[23][4]=16'h0006,loc[23][5]=16'h0004,loc[23][6]=16'hfff3,loc[23][7]=16'h0003,loc[23][8]=16'hfffe,loc[23][9]=16'hfffe,loc[23][10]=16'hfffc,loc[24][1]=16'hffff,loc[24][2]=16'hfffb,loc[24][3]=16'hfffc,loc[24][4]=16'h0001,loc[24][5]=16'h0001,loc[24][6]=16'hfffe,loc[24][7]=16'hfffe,loc[24][8]=16'h0004,loc[24][9]=16'h0000,loc[24][10]=16'h0007,loc[25][1]=16'h0004,loc[25][2]=16'h0003,loc[25][3]=16'h0005,loc[25][4]=16'h0009,loc[25][5]=16'h0002,loc[25][6]=16'hfff6,loc[25][7]=16'hfff8,loc[25][8]=16'hfff7,loc[25][9]=16'h000d,loc[25][10]=16'hfff7,loc[26][1]=16'hfffd,loc[26][2]=16'hffff,loc[26][3]=16'hfff7,loc[26][4]=16'hfffc,loc[26][5]=16'hfff3,loc[26][6]=16'hfffd,loc[26][7]=16'h000c,loc[26][8]=16'h0011,loc[26][9]=16'h0003,loc[26][10]=16'hfffd,loc[27][1]=16'h0000,loc[27][2]=16'h0004,loc[27][3]=16'h0000,loc[27][4]=16'h0009,loc[27][5]=16'h000c,loc[27][6]=16'hfff8,loc[27][7]=16'hfffe,loc[27][8]=16'hfffa,loc[27][9]=16'hfff2,loc[27][10]=16'h0007,loc[28][1]=16'h0005,loc[28][2]=16'h0004,loc[28][3]=16'hfff1,loc[28][4]=16'h0002,loc[28][5]=16'h0005,loc[28][6]=16'h0004,loc[28][7]=16'hfff4,loc[28][8]=16'h0008,loc[28][9]=16'h0009,loc[28][10]=16'hfffa,loc[29][1]=16'hffff,loc[29][2]=16'hfff8,loc[29][3]=16'h0010,loc[29][4]=16'h0013,loc[29][5]=16'hfff8,loc[29][6]=16'hfffd,loc[29][7]=16'h000a,loc[29][8]=16'h0019,loc[29][9]=16'hffe1,loc[29][10]=16'hffe7,loc[30][1]=16'hfffe,loc[30][2]=16'hfffe,loc[30][3]=16'h0006,loc[30][4]=16'h0007,loc[30][5]=16'h0007,loc[30][6]=16'hfffe,loc[30][7]=16'h0001,loc[30][8]=16'hfffb,loc[30][9]=16'hfff7,loc[30][10]=16'h0000,loc[31][1]=16'h0007,loc[31][2]=16'hffff,loc[31][3]=16'h000c,loc[31][4]=16'hfffd,loc[31][5]=16'h0005,loc[31][6]=16'h0006,loc[31][7]=16'hfff9,loc[31][8]=16'hfffb,loc[31][9]=16'hfff5,loc[31][10]=16'hfffb,loc[32][1]=16'hfffd,loc[32][2]=16'h0003,loc[32][3]=16'h0004,loc[32][4]=16'h0008,loc[32][5]=16'h0001,loc[32][6]=16'h0008,loc[32][7]=16'hffff,loc[32][8]=16'hfff2,loc[32][9]=16'h0000,loc[32][10]=16'hfffe,loc[33][1]=16'hfffa,loc[33][2]=16'hfffa,loc[33][3]=16'h0007,loc[33][4]=16'h000b,loc[33][5]=16'hffff,loc[33][6]=16'hffee,loc[33][7]=16'h000a,loc[33][8]=16'h0001,loc[33][9]=16'hffee,loc[33][10]=16'h0019,loc[34][1]=16'h000c,loc[34][2]=16'hffff,loc[34][3]=16'hfffa,loc[34][4]=16'hfff2,loc[34][5]=16'hfff6,loc[34][6]=16'h000b,loc[34][7]=16'h0005,loc[34][8]=16'hfff9,loc[34][9]=16'h0002,loc[34][10]=16'h000c,loc[35][1]=16'hfff7,loc[35][2]=16'h0007,loc[35][3]=16'h000c,loc[35][4]=16'hfffe,loc[35][5]=16'hfff9,loc[35][6]=16'hfffb,loc[35][7]=16'h0006,loc[35][8]=16'h0005,loc[35][9]=16'hffe7,loc[35][10]=16'h0015,loc[36][1]=16'hfffc,loc[36][2]=16'h0002,loc[36][3]=16'hfffe,loc[36][4]=16'hffff,loc[36][5]=16'h0009,loc[36][6]=16'h000a,loc[36][7]=16'h0001,loc[36][8]=16'hfffa,loc[36][9]=16'hfffa,loc[36][10]=16'hfffe,loc[37][1]=16'h0003,loc[37][2]=16'hfffb,loc[37][3]=16'hfffe,loc[37][4]=16'h000c,loc[37][5]=16'h0002,loc[37][6]=16'h0004,loc[37][7]=16'hfffd,loc[37][8]=16'hfff9,loc[37][9]=16'h0008,loc[37][10]=16'hfff5,loc[38][1]=16'hffff,loc[38][2]=16'hfffd,loc[38][3]=16'h0002,loc[38][4]=16'h0006,loc[38][5]=16'h0001,loc[38][6]=16'hfffe,loc[38][7]=16'hfffd,loc[38][8]=16'h0007,loc[38][9]=16'h0001,loc[38][10]=16'hfff8,loc[39][1]=16'hfffe,loc[39][2]=16'hfffd,loc[39][3]=16'hffea,loc[39][4]=16'h0010,loc[39][5]=16'hfffe,loc[39][6]=16'hfff0,loc[39][7]=16'h0000,loc[39][8]=16'h000f,loc[39][9]=16'h0017,loc[39][10]=16'hfff8,loc[40][1]=16'hfffe,loc[40][2]=16'hfff4,loc[40][3]=16'h0005,loc[40][4]=16'h000c,loc[40][5]=16'h0005,loc[40][6]=16'hfffa,loc[40][7]=16'hfffc,loc[40][8]=16'h0004,loc[40][9]=16'h0009,loc[40][10]=16'hfff6,loc[41][1]=16'h0001,loc[41][2]=16'h0008,loc[41][3]=16'h0003,loc[41][4]=16'hfff6,loc[41][5]=16'hfff8,loc[41][6]=16'h000b,loc[41][7]=16'h0003,loc[41][8]=16'hfffc,loc[41][9]=16'hfff8,loc[41][10]=16'hffff,loc[42][1]=16'h0001,loc[42][2]=16'hfffc,loc[42][3]=16'h0001,loc[42][4]=16'hfffc,loc[42][5]=16'h0006,loc[42][6]=16'hfff9,loc[42][7]=16'h0000,loc[42][8]=16'h0001,loc[42][9]=16'hfff9,loc[42][10]=16'h0009,loc[43][1]=16'h0001,loc[43][2]=16'hffff,loc[43][3]=16'h0002,loc[43][4]=16'h0000,loc[43][5]=16'h0003,loc[43][6]=16'hfffd,loc[43][7]=16'h0001,loc[43][8]=16'hffff,loc[43][9]=16'hfff6,loc[43][10]=16'h0008,loc[44][1]=16'hfff3,loc[44][2]=16'hfff8,loc[44][3]=16'h0001,loc[44][4]=16'hfff3,loc[44][5]=16'h0003,loc[44][6]=16'h0008,loc[44][7]=16'h0009,loc[44][8]=16'hffff,loc[44][9]=16'hfff1,loc[44][10]=16'h0020,loc[45][1]=16'hfffb,loc[45][2]=16'hfff4,loc[45][3]=16'hfff1,loc[45][4]=16'h0003,loc[45][5]=16'h000b,loc[45][6]=16'h0000,loc[45][7]=16'h0001,loc[45][8]=16'hfff8,loc[45][9]=16'h0016,loc[45][10]=16'h0007,loc[46][1]=16'h0000,loc[46][2]=16'h000b,loc[46][3]=16'h000c,loc[46][4]=16'hffff,loc[46][5]=16'hfff3,loc[46][6]=16'h0004,loc[46][7]=16'h0004,loc[46][8]=16'h0000,loc[46][9]=16'hfff5,loc[46][10]=16'hfffa,loc[47][1]=16'h0004,loc[47][2]=16'hfffc,loc[47][3]=16'hfffc,loc[47][4]=16'hffff,loc[47][5]=16'h0007,loc[47][6]=16'hfffc,loc[47][7]=16'hfffe,loc[47][8]=16'hfffe,loc[47][9]=16'h000b,loc[47][10]=16'h0008,loc[48][1]=16'h0003,loc[48][2]=16'h0000,loc[48][3]=16'hfffb,loc[48][4]=16'hfff8,loc[48][5]=16'hfffb,loc[48][6]=16'hfff7,loc[48][7]=16'h0003,loc[48][8]=16'h000d,loc[48][9]=16'h0000,loc[48][10]=16'h0009,loc[49][1]=16'h0003,loc[49][2]=16'hfffd,loc[49][3]=16'hfff7,loc[49][4]=16'h0009,loc[49][5]=16'h0014,loc[49][6]=16'h0004,loc[49][7]=16'hfff9,loc[49][8]=16'hfffe,loc[49][9]=16'h0006,loc[49][10]=16'hffed,loc[50][1]=16'h0012,loc[50][2]=16'h000a,loc[50][3]=16'hfffb,loc[50][4]=16'hffff,loc[50][5]=16'hfff7,loc[50][6]=16'h0000,loc[50][7]=16'hfff9,loc[50][8]=16'hfff7,loc[50][9]=16'h0009,loc[50][10]=16'hfffb,loc[51][1]=16'h0005,loc[51][2]=16'h000d,loc[51][3]=16'hfffa,loc[51][4]=16'hfff3,loc[51][5]=16'hfff6,loc[51][6]=16'h0013,loc[51][7]=16'h000d,loc[51][8]=16'hffec,loc[51][9]=16'hfff4,loc[51][10]=16'h000b,loc[52][1]=16'h0004,loc[52][2]=16'hffd9,loc[52][3]=16'hffec,loc[52][4]=16'hffad,loc[52][5]=16'hffee,loc[52][6]=16'h0043,loc[52][7]=16'h002c,loc[52][8]=16'h000e,loc[52][9]=16'h0074,loc[52][10]=16'hfff7,loc[53][1]=16'hfffd,loc[53][2]=16'h0000,loc[53][3]=16'hfffc,loc[53][4]=16'h0009,loc[53][5]=16'h0000,loc[53][6]=16'hfffd,loc[53][7]=16'h0006,loc[53][8]=16'hfff9,loc[53][9]=16'h0000,loc[53][10]=16'h0001,loc[54][1]=16'h0001,loc[54][2]=16'h0007,loc[54][3]=16'h0005,loc[54][4]=16'hfff4,loc[54][5]=16'hffff,loc[54][6]=16'h0003,loc[54][7]=16'h0004,loc[54][8]=16'hfff2,loc[54][9]=16'h0008,loc[54][10]=16'h0003,loc[55][1]=16'hfff6,loc[55][2]=16'hfff4,loc[55][3]=16'h0004,loc[55][4]=16'h0001,loc[55][5]=16'h0009,loc[55][6]=16'hfff8,loc[55][7]=16'h000a,loc[55][8]=16'h0007,loc[55][9]=16'hfff1,loc[55][10]=16'h000c,loc[56][1]=16'h0004,loc[56][2]=16'h0005,loc[56][3]=16'hfffd,loc[56][4]=16'h0008,loc[56][5]=16'hffff,loc[56][6]=16'h0002,loc[56][7]=16'hfffe,loc[56][8]=16'hfff9,loc[56][9]=16'hfffe,loc[56][10]=16'hfffc,loc[57][1]=16'h0008,loc[57][2]=16'hffff,loc[57][3]=16'h0000,loc[57][4]=16'h0015,loc[57][5]=16'hfff8,loc[57][6]=16'hfff1,loc[57][7]=16'hfff8,loc[57][8]=16'h000f,loc[57][9]=16'h0002,loc[57][10]=16'hfff3,loc[58][1]=16'hfffa,loc[58][2]=16'h0009,loc[58][3]=16'hffff,loc[58][4]=16'h0000,loc[58][5]=16'hfffb,loc[58][6]=16'hfffe,loc[58][7]=16'h000c,loc[58][8]=16'h0006,loc[58][9]=16'hfffd,loc[58][10]=16'hfff9,loc[59][1]=16'h0004,loc[59][2]=16'hfffe,loc[59][3]=16'h0008,loc[59][4]=16'h0004,loc[59][5]=16'h000e,loc[59][6]=16'hfffc,loc[59][7]=16'hfffa,loc[59][8]=16'hfffb,loc[59][9]=16'hfffd,loc[59][10]=16'hfff6,loc[60][1]=16'h0000,loc[60][2]=16'h0007,loc[60][3]=16'h0007,loc[60][4]=16'h0008,loc[60][5]=16'h0008,loc[60][6]=16'hfffb,loc[60][7]=16'hfffd,loc[60][8]=16'hfffa,loc[60][9]=16'hfff6,loc[60][10]=16'h0001,loc[61][1]=16'hfffe,loc[61][2]=16'hfffa,loc[61][3]=16'h000e,loc[61][4]=16'hfff5,loc[61][5]=16'h0012,loc[61][6]=16'h0002,loc[61][7]=16'hfff1,loc[61][8]=16'h0006,loc[61][9]=16'hfffb,loc[61][10]=16'h0003,loc[62][1]=16'h0004,loc[62][2]=16'h0008,loc[62][3]=16'h0000,loc[62][4]=16'hfff9,loc[62][5]=16'hfff9,loc[62][6]=16'h000d,loc[62][7]=16'hfff9,loc[62][8]=16'h0005,loc[62][9]=16'hfff9,loc[62][10]=16'h0001,loc[63][1]=16'hfffd,loc[63][2]=16'h0006,loc[63][3]=16'hfff9,loc[63][4]=16'hfff5,loc[63][5]=16'hfffa,loc[63][6]=16'h0001,loc[63][7]=16'hfffe,loc[63][8]=16'h000a,loc[63][9]=16'h0007,loc[63][10]=16'h0008,loc[64][1]=16'h0000,loc[64][2]=16'h0015,loc[64][3]=16'h0001,loc[64][4]=16'h0001,loc[64][5]=16'hffee,loc[64][6]=16'h0004,loc[64][7]=16'hfffc,loc[64][8]=16'h0003,loc[64][9]=16'h0009,loc[64][10]=16'hfff8,loc[65][1]=16'hffff,loc[65][2]=16'h0010,loc[65][3]=16'hfff7,loc[65][4]=16'hfffa,loc[65][5]=16'hfffd,loc[65][6]=16'h000e,loc[65][7]=16'h0001,loc[65][8]=16'h0003,loc[65][9]=16'h0003,loc[65][10]=16'hfff2,loc[66][1]=16'h0002,loc[66][2]=16'hffff,loc[66][3]=16'hfffc,loc[66][4]=16'h0008,loc[66][5]=16'hfffd,loc[66][6]=16'hfff8,loc[66][7]=16'h0001,loc[66][8]=16'h0004,loc[66][9]=16'h0007,loc[66][10]=16'hfffe,loc[67][1]=16'h000b,loc[67][2]=16'h0002,loc[67][3]=16'hfffb,loc[67][4]=16'h0009,loc[67][5]=16'h0003,loc[67][6]=16'hfff9,loc[67][7]=16'hfff6,loc[67][8]=16'hfffe,loc[67][9]=16'hfffb,loc[67][10]=16'hfffe,loc[68][1]=16'h0003,loc[68][2]=16'h0007,loc[68][3]=16'h0006,loc[68][4]=16'h0007,loc[68][5]=16'hfffc,loc[68][6]=16'hfffc,loc[68][7]=16'hfffb,loc[68][8]=16'h0009,loc[68][9]=16'hfff4,loc[68][10]=16'hfffa,loc[69][1]=16'h0005,loc[69][2]=16'hfffd,loc[69][3]=16'hfff8,loc[69][4]=16'h0002,loc[69][5]=16'h0001,loc[69][6]=16'hfff9,loc[69][7]=16'h0000,loc[69][8]=16'h0008,loc[69][9]=16'h0006,loc[69][10]=16'hffff,loc[70][1]=16'h000e,loc[70][2]=16'h0005,loc[70][3]=16'h0007,loc[70][4]=16'hfffc,loc[70][5]=16'hfff8,loc[70][6]=16'h0007,loc[70][7]=16'hfffb,loc[70][8]=16'hfff2,loc[70][9]=16'h0005,loc[70][10]=16'hfffe,loc[71][1]=16'hfffd,loc[71][2]=16'h0002,loc[71][3]=16'h0003,loc[71][4]=16'hfff8,loc[71][5]=16'h0002,loc[71][6]=16'h0001,loc[71][7]=16'h0002,loc[71][8]=16'hfffb,loc[71][9]=16'hfffa,loc[71][10]=16'h0009,loc[72][1]=16'h0003,loc[72][2]=16'hffff,loc[72][3]=16'h0002,loc[72][4]=16'hfffa,loc[72][5]=16'hffff,loc[72][6]=16'h0007,loc[72][7]=16'hfffa,loc[72][8]=16'h0005,loc[72][9]=16'h0004,loc[72][10]=16'hfffa,loc[73][1]=16'h0000,loc[73][2]=16'hfffb,loc[73][3]=16'h0001,loc[73][4]=16'hffff,loc[73][5]=16'h0001,loc[73][6]=16'h0000,loc[73][7]=16'h0001,loc[73][8]=16'h0001,loc[73][9]=16'hfffc,loc[73][10]=16'h0001,loc[74][1]=16'h0003,loc[74][2]=16'hffff,loc[74][3]=16'hfffe,loc[74][4]=16'h0003,loc[74][5]=16'hfff6,loc[74][6]=16'hfffd,loc[74][7]=16'h000e,loc[74][8]=16'h0000,loc[74][9]=16'hfffb,loc[74][10]=16'h0004,loc[75][1]=16'h0003,loc[75][2]=16'h0000,loc[75][3]=16'h0001,loc[75][4]=16'h0007,loc[75][5]=16'hfffb,loc[75][6]=16'hfff9,loc[75][7]=16'h0004,loc[75][8]=16'h0000,loc[75][9]=16'hfff6,loc[75][10]=16'h0004,loc[76][1]=16'hfffe,loc[76][2]=16'hfffc,loc[76][3]=16'h0002,loc[76][4]=16'hfff9,loc[76][5]=16'hfffc,loc[76][6]=16'hfffb,loc[76][7]=16'hfff7,loc[76][8]=16'h000c,loc[76][9]=16'h000e,loc[76][10]=16'hffff,loc[77][1]=16'h0003,loc[77][2]=16'hfff8,loc[77][3]=16'hfffb,loc[77][4]=16'h0005,loc[77][5]=16'h0002,loc[77][6]=16'h0000,loc[77][7]=16'h0000,loc[77][8]=16'h0005,loc[77][9]=16'hfffd,loc[77][10]=16'h0003,loc[78][1]=16'h0006,loc[78][2]=16'h0001,loc[78][3]=16'hfff4,loc[78][4]=16'hfffb,loc[78][5]=16'hfffc,loc[78][6]=16'h000a,loc[78][7]=16'hfff8,loc[78][8]=16'h0011,loc[78][9]=16'hffeb,loc[78][10]=16'h000e,loc[79][1]=16'hffff,loc[79][2]=16'h0007,loc[79][3]=16'h0005,loc[79][4]=16'h0005,loc[79][5]=16'hfff9,loc[79][6]=16'hfffa,loc[79][7]=16'h0007,loc[79][8]=16'h0000,loc[79][9]=16'hfff9,loc[79][10]=16'h0000,loc[80][1]=16'h0001,loc[80][2]=16'h0000,loc[80][3]=16'h0013,loc[80][4]=16'h0002,loc[80][5]=16'h0000,loc[80][6]=16'h0001,loc[80][7]=16'h0001,loc[80][8]=16'hfffd,loc[80][9]=16'hfff6,loc[80][10]=16'hfffc,loc[81][1]=16'h0004,loc[81][2]=16'hfffa,loc[81][3]=16'h0000,loc[81][4]=16'hfff7,loc[81][5]=16'h0004,loc[81][6]=16'h0000,loc[81][7]=16'hfff8,loc[81][8]=16'h0008,loc[81][9]=16'h0001,loc[81][10]=16'h0009,loc[82][1]=16'hfffd,loc[82][2]=16'h0007,loc[82][3]=16'h0005,loc[82][4]=16'hfffa,loc[82][5]=16'h0000,loc[82][6]=16'h0006,loc[82][7]=16'hfff4,loc[82][8]=16'h0001,loc[82][9]=16'h0004,loc[82][10]=16'hfffd,loc[83][1]=16'h0004,loc[83][2]=16'h000a,loc[83][3]=16'h0002,loc[83][4]=16'hfffe,loc[83][5]=16'hfff9,loc[83][6]=16'hffff,loc[83][7]=16'hfffd,loc[83][8]=16'h0002,loc[83][9]=16'h0001,loc[83][10]=16'hfffb,loc[84][1]=16'h0001,loc[84][2]=16'hfffc,loc[84][3]=16'h0004,loc[84][4]=16'h0005,loc[84][5]=16'h0005,loc[84][6]=16'h0002,loc[84][7]=16'hfffc,loc[84][8]=16'hfffb,loc[84][9]=16'hfffe,loc[84][10]=16'hfff8,loc[85][1]=16'hfffd,loc[85][2]=16'h0002,loc[85][3]=16'hfffb,loc[85][4]=16'h0000,loc[85][5]=16'h0000,loc[85][6]=16'hffff,loc[85][7]=16'h0002,loc[85][8]=16'hfffe,loc[85][9]=16'h000a,loc[85][10]=16'hffff,loc[86][1]=16'hfffe,loc[86][2]=16'h0002,loc[86][3]=16'hfffd,loc[86][4]=16'h0005,loc[86][5]=16'h0008,loc[86][6]=16'h0005,loc[86][7]=16'hfffd,loc[86][8]=16'hfffa,loc[86][9]=16'hfffa,loc[86][10]=16'hfffd,loc[87][1]=16'h000a,loc[87][2]=16'hfffb,loc[87][3]=16'hfffe,loc[87][4]=16'h0007,loc[87][5]=16'hfff7,loc[87][6]=16'h000f,loc[87][7]=16'h0005,loc[87][8]=16'h0006,loc[87][9]=16'hfff4,loc[87][10]=16'hfff3,loc[88][1]=16'h0004,loc[88][2]=16'h0008,loc[88][3]=16'hfffc,loc[88][4]=16'h000b,loc[88][5]=16'hfffe,loc[88][6]=16'hfffb,loc[88][7]=16'h0002,loc[88][8]=16'hfff4,loc[88][9]=16'h0000,loc[88][10]=16'h0002,loc[89][1]=16'h0005,loc[89][2]=16'hfffd,loc[89][3]=16'hfffd,loc[89][4]=16'hfff4,loc[89][5]=16'h0006,loc[89][6]=16'h0002,loc[89][7]=16'hfffe,loc[89][8]=16'h000b,loc[89][9]=16'h0005,loc[89][10]=16'hfffa,loc[90][1]=16'hfffd,loc[90][2]=16'hfffe,loc[90][3]=16'hfffc,loc[90][4]=16'hfff5,loc[90][5]=16'h0001,loc[90][6]=16'h0008,loc[90][7]=16'h0011,loc[90][8]=16'hfffd,loc[90][9]=16'hffff,loc[90][10]=16'hfffe,loc[91][1]=16'h0007,loc[91][2]=16'h0005,loc[91][3]=16'h0003,loc[91][4]=16'hfff5,loc[91][5]=16'hfffc,loc[91][6]=16'h0001,loc[91][7]=16'h0000,loc[91][8]=16'h0005,loc[91][9]=16'hfff8,loc[91][10]=16'h0003,loc[92][1]=16'hffff,loc[92][2]=16'h0001,loc[92][3]=16'hfff8,loc[92][4]=16'h0007,loc[92][5]=16'hffff,loc[92][6]=16'h0002,loc[92][7]=16'h0003,loc[92][8]=16'hfffc,loc[92][9]=16'hfffe,loc[92][10]=16'h0004,loc[93][1]=16'hfffe,loc[93][2]=16'hfffc,loc[93][3]=16'h0004,loc[93][4]=16'h0009,loc[93][5]=16'hfff7,loc[93][6]=16'h0003,loc[93][7]=16'hffff,loc[93][8]=16'h0005,loc[93][9]=16'h0001,loc[93][10]=16'hfffc,loc[94][1]=16'h0005,loc[94][2]=16'hfffd,loc[94][3]=16'hfffb,loc[94][4]=16'hfffe,loc[94][5]=16'hfffa,loc[94][6]=16'h000a,loc[94][7]=16'h0005,loc[94][8]=16'h0009,loc[94][9]=16'hfff9,loc[94][10]=16'hfffc,loc[95][1]=16'hffff,loc[95][2]=16'hffef,loc[95][3]=16'hffe8,loc[95][4]=16'h0014,loc[95][5]=16'h0005,loc[95][6]=16'h0006,loc[95][7]=16'hfffd,loc[95][8]=16'h0009,loc[95][9]=16'hfffc,loc[95][10]=16'h0002,loc[96][1]=16'hffff,loc[96][2]=16'hfff9,loc[96][3]=16'h000a,loc[96][4]=16'hfff6,loc[96][5]=16'hfffd,loc[96][6]=16'h0003,loc[96][7]=16'h0004,loc[96][8]=16'h0007,loc[96][9]=16'hfff5,loc[96][10]=16'h0008,loc[97][1]=16'h0000,loc[97][2]=16'h0007,loc[97][3]=16'hffff,loc[97][4]=16'h0002,loc[97][5]=16'hfffd,loc[97][6]=16'hfffc,loc[97][7]=16'hfffc,loc[97][8]=16'hfffb,loc[97][9]=16'h0004,loc[97][10]=16'h0004,loc[98][1]=16'h0009,loc[98][2]=16'hffff,loc[98][3]=16'hfff6,loc[98][4]=16'h0006,loc[98][5]=16'h0004,loc[98][6]=16'hfff5,loc[98][7]=16'h000a,loc[98][8]=16'h0008,loc[98][9]=16'hfff0,loc[98][10]=16'h0005,loc[99][1]=16'h0003,loc[99][2]=16'h0002,loc[99][3]=16'hfff8,loc[99][4]=16'hfffb,loc[99][5]=16'hfff7,loc[99][6]=16'h0001,loc[99][7]=16'h0006,loc[99][8]=16'h0004,loc[99][9]=16'h0007,loc[99][10]=16'h0000,loc[100][1]=16'h0000,loc[100][2]=16'h0006,loc[100][3]=16'h0008,loc[100][4]=16'hfffd,loc[100][5]=16'h0004,loc[100][6]=16'h0003,loc[100][7]=16'hfff8,loc[100][8]=16'hfff5,loc[100][9]=16'h0003,loc[100][10]=16'hffff,loc[101][1]=16'hfffb,loc[101][2]=16'h0006,loc[101][3]=16'h0006,loc[101][4]=16'hfffd,loc[101][5]=16'h0006,loc[101][6]=16'hfffc,loc[101][7]=16'h0008,loc[101][8]=16'hfffc,loc[101][9]=16'hfffc,loc[101][10]=16'hfffd,loc[102][1]=16'hfffe,loc[102][2]=16'hfff6,loc[102][3]=16'hffff,loc[102][4]=16'h0007,loc[102][5]=16'hfffe,loc[102][6]=16'h0000,loc[102][7]=16'h000a,loc[102][8]=16'h0005,loc[102][9]=16'h0002,loc[102][10]=16'hfff9,loc[103][1]=16'h000e,loc[103][2]=16'h0001,loc[103][3]=16'hfff9,loc[103][4]=16'h000c,loc[103][5]=16'hffea,loc[103][6]=16'h0005,loc[103][7]=16'h0006,loc[103][8]=16'hffef,loc[103][9]=16'h0014,loc[103][10]=16'hffff,loc[104][1]=16'h0002,loc[104][2]=16'h0001,loc[104][3]=16'hfff9,loc[104][4]=16'hffff,loc[104][5]=16'hfffc,loc[104][6]=16'h0008,loc[104][7]=16'h0001,loc[104][8]=16'hfffc,loc[104][9]=16'h0007,loc[104][10]=16'hfffd,loc[105][1]=16'hfff8,loc[105][2]=16'hfff7,loc[105][3]=16'h000c,loc[105][4]=16'h0007,loc[105][5]=16'hfffc,loc[105][6]=16'h0013,loc[105][7]=16'h0002,loc[105][8]=16'hffee,loc[105][9]=16'h0016,loc[105][10]=16'hffe5,loc[106][1]=16'h0001,loc[106][2]=16'h0000,loc[106][3]=16'hffff,loc[106][4]=16'hfff8,loc[106][5]=16'hfffb,loc[106][6]=16'hfffe,loc[106][7]=16'hfff3,loc[106][8]=16'h000c,loc[106][9]=16'h0020,loc[106][10]=16'hfff5,loc[107][1]=16'hfffd,loc[107][2]=16'h0004,loc[107][3]=16'h0004,loc[107][4]=16'hfffd,loc[107][5]=16'hfffa,loc[107][6]=16'h000b,loc[107][7]=16'h0000,loc[107][8]=16'hfffd,loc[107][9]=16'h0000,loc[107][10]=16'h0000,loc[108][1]=16'h0002,loc[108][2]=16'hfffd,loc[108][3]=16'h0009,loc[108][4]=16'hfffe,loc[108][5]=16'hfffd,loc[108][6]=16'h000b,loc[108][7]=16'hfffc,loc[108][8]=16'h000e,loc[108][9]=16'hfffe,loc[108][10]=16'hfff3,loc[109][1]=16'h0000,loc[109][2]=16'hfff8,loc[109][3]=16'hfffb,loc[109][4]=16'h0005,loc[109][5]=16'h0000,loc[109][6]=16'h0000,loc[109][7]=16'h0006,loc[109][8]=16'h0009,loc[109][9]=16'h0006,loc[109][10]=16'hfff6,loc[110][1]=16'h0008,loc[110][2]=16'hffff,loc[110][3]=16'hfffb,loc[110][4]=16'hfff2,loc[110][5]=16'hfffd,loc[110][6]=16'h0003,loc[110][7]=16'h0000,loc[110][8]=16'h000b,loc[110][9]=16'hfffd,loc[110][10]=16'h0005,loc[111][1]=16'h0000,loc[111][2]=16'h0005,loc[111][3]=16'hffff,loc[111][4]=16'hffff,loc[111][5]=16'h0002,loc[111][6]=16'h0008,loc[111][7]=16'hfffc,loc[111][8]=16'h0007,loc[111][9]=16'hfff0,loc[111][10]=16'hfffe,loc[112][1]=16'hfffc,loc[112][2]=16'hfff9,loc[112][3]=16'h0004,loc[112][4]=16'hffff,loc[112][5]=16'hfffe,loc[112][6]=16'hfffa,loc[112][7]=16'h000a,loc[112][8]=16'h0008,loc[112][9]=16'hfff9,loc[112][10]=16'h0006,loc[113][1]=16'h0004,loc[113][2]=16'hfff9,loc[113][3]=16'h000a,loc[113][4]=16'h0009,loc[113][5]=16'hfffa,loc[113][6]=16'hfffe,loc[113][7]=16'h0006,loc[113][8]=16'h0006,loc[113][9]=16'hfff7,loc[113][10]=16'hfff5,loc[114][1]=16'h0004,loc[114][2]=16'hffff,loc[114][3]=16'hfff9,loc[114][4]=16'h0002,loc[114][5]=16'hfffa,loc[114][6]=16'hffff,loc[114][7]=16'h0009,loc[114][8]=16'h0004,loc[114][9]=16'hffff,loc[114][10]=16'h0002,loc[115][1]=16'h0002,loc[115][2]=16'hfff8,loc[115][3]=16'hfffe,loc[115][4]=16'h0003,loc[115][5]=16'h0004,loc[115][6]=16'hfffb,loc[115][7]=16'h0008,loc[115][8]=16'hfffd,loc[115][9]=16'hfff8,loc[115][10]=16'h000b,loc[116][1]=16'h0002,loc[116][2]=16'h0004,loc[116][3]=16'h0004,loc[116][4]=16'hfffe,loc[116][5]=16'hfffa,loc[116][6]=16'hfffb,loc[116][7]=16'hfffe,loc[116][8]=16'h0001,loc[116][9]=16'h0000,loc[116][10]=16'h0002,loc[117][1]=16'h002a,loc[117][2]=16'h000d,loc[117][3]=16'h000f,loc[117][4]=16'hffe9,loc[117][5]=16'hffe1,loc[117][6]=16'hfff1,loc[117][7]=16'h001c,loc[117][8]=16'hffcd,loc[117][9]=16'hffce,loc[117][10]=16'h004a,loc[118][1]=16'h0002,loc[118][2]=16'h0001,loc[118][3]=16'hfff8,loc[118][4]=16'hffff,loc[118][5]=16'hfffd,loc[118][6]=16'hffff,loc[118][7]=16'h0005,loc[118][8]=16'h0000,loc[118][9]=16'h0005,loc[118][10]=16'hffff,loc[119][1]=16'h0001,loc[119][2]=16'h0003,loc[119][3]=16'hfff6,loc[119][4]=16'hfffc,loc[119][5]=16'hfffd,loc[119][6]=16'hfffe,loc[119][7]=16'h0006,loc[119][8]=16'h0001,loc[119][9]=16'hfff6,loc[119][10]=16'h0010,loc[120][1]=16'h0006,loc[120][2]=16'h0002,loc[120][3]=16'hfffc,loc[120][4]=16'hfffe,loc[120][5]=16'hfff7,loc[120][6]=16'h0002,loc[120][7]=16'hfff9,loc[120][8]=16'h0002,loc[120][9]=16'h0002,loc[120][10]=16'h0007,loc[121][1]=16'h0001,loc[121][2]=16'hfff7,loc[121][3]=16'hfffa,loc[121][4]=16'hfffa,loc[121][5]=16'hfff9,loc[121][6]=16'hffff,loc[121][7]=16'h0002,loc[121][8]=16'h0007,loc[121][9]=16'h0003,loc[121][10]=16'h0012,loc[122][1]=16'h0003,loc[122][2]=16'h0003,loc[122][3]=16'hffff,loc[122][4]=16'h0001,loc[122][5]=16'h000d,loc[122][6]=16'h0009,loc[122][7]=16'hfff7,loc[122][8]=16'hfffa,loc[122][9]=16'hfff6,loc[122][10]=16'h0000,loc[123][1]=16'hfff7,loc[123][2]=16'hfffc,loc[123][3]=16'h0009,loc[123][4]=16'h0008,loc[123][5]=16'h0007,loc[123][6]=16'hfff9,loc[123][7]=16'hfff8,loc[123][8]=16'h0002,loc[123][9]=16'h0001,loc[123][10]=16'h0004,loc[124][1]=16'h0003,loc[124][2]=16'h0002,loc[124][3]=16'hfffb,loc[124][4]=16'h0005,loc[124][5]=16'hfff9,loc[124][6]=16'h0000,loc[124][7]=16'h0003,loc[124][8]=16'h0007,loc[124][9]=16'hfffa,loc[124][10]=16'h0000,loc[125][1]=16'h0001,loc[125][2]=16'h0003,loc[125][3]=16'h0006,loc[125][4]=16'h0005,loc[125][5]=16'hfffe,loc[125][6]=16'hfffc,loc[125][7]=16'hfffa,loc[125][8]=16'hfff7,loc[125][9]=16'h0006,loc[125][10]=16'h0002,loc[126][1]=16'h0000,loc[126][2]=16'h0004,loc[126][3]=16'hfffc,loc[126][4]=16'h0002,loc[126][5]=16'hfff9,loc[126][6]=16'hfffa,loc[126][7]=16'h0001,loc[126][8]=16'h0001,loc[126][9]=16'h0001,loc[126][10]=16'h0009,loc[127][1]=16'hfff9,loc[127][2]=16'hfff9,loc[127][3]=16'h0001,loc[127][4]=16'h0001,loc[127][5]=16'hffff,loc[127][6]=16'hfffe,loc[127][7]=16'h0005,loc[127][8]=16'h0005,loc[127][9]=16'h0002,loc[127][10]=16'h0000,loc[128][1]=16'h001d,loc[128][2]=16'h0019,loc[128][3]=16'h0008,loc[128][4]=16'hffef,loc[128][5]=16'hffe2,loc[128][6]=16'h0010,loc[128][7]=16'hffd8,loc[128][8]=16'h0002,loc[128][9]=16'h0008,loc[128][10]=16'h001b,loc[129][1]=16'hfffb,loc[129][2]=16'h0002,loc[129][3]=16'h0008,loc[129][4]=16'h0003,loc[129][5]=16'h0000,loc[129][6]=16'hfffc,loc[129][7]=16'h0006,loc[129][8]=16'hfffd,loc[129][9]=16'hfffc,loc[129][10]=16'hfffc,loc[130][1]=16'h0006,loc[130][2]=16'hfffd,loc[130][3]=16'hfffb,loc[130][4]=16'h0006,loc[130][5]=16'h0004,loc[130][6]=16'hfff5,loc[130][7]=16'h0001,loc[130][8]=16'hfffe,loc[130][9]=16'h0004,loc[130][10]=16'h0001,loc[131][1]=16'h0006,loc[131][2]=16'h0003,loc[131][3]=16'h0000,loc[131][4]=16'h0003,loc[131][5]=16'h0009,loc[131][6]=16'h000a,loc[131][7]=16'hfff6,loc[131][8]=16'hfffa,loc[131][9]=16'hfffa,loc[131][10]=16'hfffa,loc[132][1]=16'h0006,loc[132][2]=16'h0003,loc[132][3]=16'h0006,loc[132][4]=16'h0008,loc[132][5]=16'hfffa,loc[132][6]=16'h0002,loc[132][7]=16'hfffd,loc[132][8]=16'hfff9,loc[132][9]=16'hfffd,loc[132][10]=16'hfffc,loc[133][1]=16'h0002,loc[133][2]=16'h0002,loc[133][3]=16'h0005,loc[133][4]=16'h0004,loc[133][5]=16'h0002,loc[133][6]=16'h0006,loc[133][7]=16'h0004,loc[133][8]=16'hffee,loc[133][9]=16'h0002,loc[133][10]=16'hfffa,loc[134][1]=16'h0008,loc[134][2]=16'h0000,loc[134][3]=16'h0000,loc[134][4]=16'h0004,loc[134][5]=16'hfffb,loc[134][6]=16'hfffa,loc[134][7]=16'h0002,loc[134][8]=16'h0000,loc[134][9]=16'hfff7,loc[134][10]=16'h0004,loc[135][1]=16'hffff,loc[135][2]=16'h000a,loc[135][3]=16'hfffd,loc[135][4]=16'hfffc,loc[135][5]=16'hfffd,loc[135][6]=16'hfff3,loc[135][7]=16'h0007,loc[135][8]=16'h0000,loc[135][9]=16'h0001,loc[135][10]=16'h0005,loc[136][1]=16'h000a,loc[136][2]=16'h0005,loc[136][3]=16'hfffb,loc[136][4]=16'hfffb,loc[136][5]=16'hfffa,loc[136][6]=16'h000f,loc[136][7]=16'hfff0,loc[136][8]=16'h0001,loc[136][9]=16'h0003,loc[136][10]=16'hfffa,loc[137][1]=16'hffff,loc[137][2]=16'h0007,loc[137][3]=16'hfff9,loc[137][4]=16'h0007,loc[137][5]=16'h0000,loc[137][6]=16'h0004,loc[137][7]=16'h0001,loc[137][8]=16'hfffc,loc[137][9]=16'hfff7,loc[137][10]=16'h0007,loc[138][1]=16'hfffa,loc[138][2]=16'hfff9,loc[138][3]=16'hffff,loc[138][4]=16'h0004,loc[138][5]=16'hfffb,loc[138][6]=16'h0005,loc[138][7]=16'h0003,loc[138][8]=16'h000c,loc[138][9]=16'hfff5,loc[138][10]=16'h0007,loc[139][1]=16'h0003,loc[139][2]=16'h0002,loc[139][3]=16'h0003,loc[139][4]=16'h0000,loc[139][5]=16'hfffd,loc[139][6]=16'hfff7,loc[139][7]=16'hfff8,loc[139][8]=16'hfffd,loc[139][9]=16'h000d,loc[139][10]=16'h0000,loc[140][1]=16'hfff9,loc[140][2]=16'hfffd,loc[140][3]=16'h0000,loc[140][4]=16'hfffe,loc[140][5]=16'h000e,loc[140][6]=16'hfff8,loc[140][7]=16'hffff,loc[140][8]=16'h0001,loc[140][9]=16'h0013,loc[140][10]=16'hfff6,loc[141][1]=16'h0003,loc[141][2]=16'h0018,loc[141][3]=16'h0000,loc[141][4]=16'h000a,loc[141][5]=16'hfff0,loc[141][6]=16'h0006,loc[141][7]=16'hffe2,loc[141][8]=16'hfff5,loc[141][9]=16'h000f,loc[141][10]=16'h000a,loc[142][1]=16'hfff6,loc[142][2]=16'h0000,loc[142][3]=16'hffff,loc[142][4]=16'hfff6,loc[142][5]=16'h0006,loc[142][6]=16'hfff9,loc[142][7]=16'hfff7,loc[142][8]=16'h0009,loc[142][9]=16'h0004,loc[142][10]=16'h0012,loc[143][1]=16'h000a,loc[143][2]=16'h005a,loc[143][3]=16'hffcc,loc[143][4]=16'hfff1,loc[143][5]=16'h000c,loc[143][6]=16'h0006,loc[143][7]=16'hffc9,loc[143][8]=16'hffe5,loc[143][9]=16'h0026,loc[143][10]=16'h0002,loc[144][1]=16'h0005,loc[144][2]=16'hfffe,loc[144][3]=16'h0009,loc[144][4]=16'hfff9,loc[144][5]=16'h0009,loc[144][6]=16'h0001,loc[144][7]=16'hffef,loc[144][8]=16'hfffd,loc[144][9]=16'h0008,loc[144][10]=16'hffff,loc[145][1]=16'h0000,loc[145][2]=16'hfffb,loc[145][3]=16'hfffa,loc[145][4]=16'h0002,loc[145][5]=16'h0002,loc[145][6]=16'hfff8,loc[145][7]=16'h0009,loc[145][8]=16'h0003,loc[145][9]=16'h0001,loc[145][10]=16'h0004,loc[146][1]=16'hffff,loc[146][2]=16'hfffe,loc[146][3]=16'hfffd,loc[146][4]=16'hfffb,loc[146][5]=16'hfff9,loc[146][6]=16'h0003,loc[146][7]=16'h0007,loc[146][8]=16'h0005,loc[146][9]=16'h0007,loc[146][10]=16'hffff,loc[147][1]=16'h0002,loc[147][2]=16'h0000,loc[147][3]=16'h0004,loc[147][4]=16'hfff7,loc[147][5]=16'hffff,loc[147][6]=16'h000d,loc[147][7]=16'h0000,loc[147][8]=16'hfffe,loc[147][9]=16'hfff9,loc[147][10]=16'h0002,loc[148][1]=16'h0004,loc[148][2]=16'h0008,loc[148][3]=16'hfffa,loc[148][4]=16'hfffc,loc[148][5]=16'hfffe,loc[148][6]=16'h0000,loc[148][7]=16'hfffe,loc[148][8]=16'h0002,loc[148][9]=16'h0004,loc[148][10]=16'h0002,loc[149][1]=16'hffff,loc[149][2]=16'h000d,loc[149][3]=16'hfffb,loc[149][4]=16'h0004,loc[149][5]=16'hfff7,loc[149][6]=16'hfffe,loc[149][7]=16'h0005,loc[149][8]=16'h0000,loc[149][9]=16'hfffc,loc[149][10]=16'h0001,loc[150][1]=16'h0003,loc[150][2]=16'h0000,loc[150][3]=16'h0002,loc[150][4]=16'hfff8,loc[150][5]=16'h0000,loc[150][6]=16'h0007,loc[150][7]=16'h0001,loc[150][8]=16'h0006,loc[150][9]=16'hffff,loc[150][10]=16'hfffa,loc[151][1]=16'hfff6,loc[151][2]=16'hffef,loc[151][3]=16'h0005,loc[151][4]=16'h0003,loc[151][5]=16'hfffc,loc[151][6]=16'hfffb,loc[151][7]=16'h0004,loc[151][8]=16'h0017,loc[151][9]=16'hfff4,loc[151][10]=16'h0006,loc[152][1]=16'h0003,loc[152][2]=16'hfff2,loc[152][3]=16'hfffd,loc[152][4]=16'h0009,loc[152][5]=16'h0002,loc[152][6]=16'hfff5,loc[152][7]=16'h0003,loc[152][8]=16'h0000,loc[152][9]=16'h0007,loc[152][10]=16'h0005,loc[153][1]=16'h0001,loc[153][2]=16'h0006,loc[153][3]=16'hfffa,loc[153][4]=16'hfffc,loc[153][5]=16'hfffe,loc[153][6]=16'h0002,loc[153][7]=16'h0002,loc[153][8]=16'h0005,loc[153][9]=16'h0002,loc[153][10]=16'hfffe,loc[154][1]=16'hfffc,loc[154][2]=16'hfff9,loc[154][3]=16'h0002,loc[154][4]=16'h0008,loc[154][5]=16'h0008,loc[154][6]=16'hfffe,loc[154][7]=16'hfffc,loc[154][8]=16'hffff,loc[154][9]=16'h0002,loc[154][10]=16'hffff,loc[155][1]=16'h0006,loc[155][2]=16'hfff9,loc[155][3]=16'h0009,loc[155][4]=16'hfffe,loc[155][5]=16'h0006,loc[155][6]=16'h0004,loc[155][7]=16'hfff7,loc[155][8]=16'h0009,loc[155][9]=16'hfff1,loc[155][10]=16'hffff,loc[156][1]=16'h0003,loc[156][2]=16'h0002,loc[156][3]=16'h0002,loc[156][4]=16'hffff,loc[156][5]=16'h0005,loc[156][6]=16'h0001,loc[156][7]=16'hfff8,loc[156][8]=16'hfffb,loc[156][9]=16'hfffc,loc[156][10]=16'h0005,loc[157][1]=16'hfffd,loc[157][2]=16'h0016,loc[157][3]=16'hfff6,loc[157][4]=16'hfff0,loc[157][5]=16'hfffd,loc[157][6]=16'h0004,loc[157][7]=16'hffff,loc[157][8]=16'h0005,loc[157][9]=16'h0005,loc[157][10]=16'h0000,loc[158][1]=16'hfff9,loc[158][2]=16'hfff7,loc[158][3]=16'hffff,loc[158][4]=16'hffff,loc[158][5]=16'h0008,loc[158][6]=16'hfffe,loc[158][7]=16'h0003,loc[158][8]=16'h0002,loc[158][9]=16'h000e,loc[158][10]=16'hfffc,loc[159][1]=16'h0003,loc[159][2]=16'h0005,loc[159][3]=16'hfff1,loc[159][4]=16'h0009,loc[159][5]=16'hfff5,loc[159][6]=16'hfffd,loc[159][7]=16'h0009,loc[159][8]=16'hffff,loc[159][9]=16'h0001,loc[159][10]=16'h0004,loc[160][1]=16'hffff,loc[160][2]=16'hfffb,loc[160][3]=16'h0004,loc[160][4]=16'h0006,loc[160][5]=16'hfffd,loc[160][6]=16'hfffe,loc[160][7]=16'hffff,loc[160][8]=16'h0001,loc[160][9]=16'h0003,loc[160][10]=16'hfffb,loc[161][1]=16'hffeb,loc[161][2]=16'hffd9,loc[161][3]=16'hfff6,loc[161][4]=16'hffe4,loc[161][5]=16'h002a,loc[161][6]=16'hffe9,loc[161][7]=16'h0005,loc[161][8]=16'h0010,loc[161][9]=16'h0019,loc[161][10]=16'h0023,loc[162][1]=16'hfff8,loc[162][2]=16'h0003,loc[162][3]=16'hfffb,loc[162][4]=16'h0001,loc[162][5]=16'hfffa,loc[162][6]=16'hfff9,loc[162][7]=16'h0008,loc[162][8]=16'hfffe,loc[162][9]=16'h0002,loc[162][10]=16'h000c,loc[163][1]=16'h000a,loc[163][2]=16'hffeb,loc[163][3]=16'h0000,loc[163][4]=16'h0004,loc[163][5]=16'h000b,loc[163][6]=16'hffeb,loc[163][7]=16'h0008,loc[163][8]=16'hfffa,loc[163][9]=16'h0002,loc[163][10]=16'h000c,loc[164][1]=16'h0003,loc[164][2]=16'h0009,loc[164][3]=16'hfffb,loc[164][4]=16'h0001,loc[164][5]=16'hfffe,loc[164][6]=16'hffff,loc[164][7]=16'h000b,loc[164][8]=16'hfff4,loc[164][9]=16'hfffa,loc[164][10]=16'h0009,loc[165][1]=16'h0001,loc[165][2]=16'h0006,loc[165][3]=16'hfffc,loc[165][4]=16'h0008,loc[165][5]=16'h0005,loc[165][6]=16'h0004,loc[165][7]=16'hffff,loc[165][8]=16'hfff9,loc[165][9]=16'h0004,loc[165][10]=16'hfff6,loc[166][1]=16'h0003,loc[166][2]=16'h0001,loc[166][3]=16'hfffb,loc[166][4]=16'h0004,loc[166][5]=16'h0002,loc[166][6]=16'h0003,loc[166][7]=16'hfffa,loc[166][8]=16'hffff,loc[166][9]=16'hfffb,loc[166][10]=16'h0004,loc[167][1]=16'h0002,loc[167][2]=16'h0002,loc[167][3]=16'hffff,loc[167][4]=16'hfffe,loc[167][5]=16'hfffe,loc[167][6]=16'hfffa,loc[167][7]=16'hffff,loc[167][8]=16'h0005,loc[167][9]=16'h0000,loc[167][10]=16'h0002,loc[168][1]=16'h0003,loc[168][2]=16'h0004,loc[168][3]=16'hfffb,loc[168][4]=16'hfff8,loc[168][5]=16'hfffb,loc[168][6]=16'hfffc,loc[168][7]=16'h0002,loc[168][8]=16'h0005,loc[168][9]=16'h0004,loc[168][10]=16'h0006,loc[169][1]=16'h0008,loc[169][2]=16'h0003,loc[169][3]=16'hfffc,loc[169][4]=16'hfff8,loc[169][5]=16'h0005,loc[169][6]=16'h0002,loc[169][7]=16'hfff5,loc[169][8]=16'h000b,loc[169][9]=16'h0006,loc[169][10]=16'hfff4,loc[170][1]=16'h0004,loc[170][2]=16'h0006,loc[170][3]=16'h0002,loc[170][4]=16'hfff7,loc[170][5]=16'h0004,loc[170][6]=16'h0002,loc[170][7]=16'hfffe,loc[170][8]=16'hffff,loc[170][9]=16'hfff2,loc[170][10]=16'h000a,loc[171][1]=16'h0000,loc[171][2]=16'h0000,loc[171][3]=16'h000d,loc[171][4]=16'hfff9,loc[171][5]=16'hfff7,loc[171][6]=16'h000b,loc[171][7]=16'h0006,loc[171][8]=16'h0005,loc[171][9]=16'h0000,loc[171][10]=16'hfff2,loc[172][1]=16'hfffd,loc[172][2]=16'hfff9,loc[172][3]=16'h000c,loc[172][4]=16'hfffa,loc[172][5]=16'h0002,loc[172][6]=16'h0005,loc[172][7]=16'hfffb,loc[172][8]=16'h0008,loc[172][9]=16'h0002,loc[172][10]=16'hfffc,loc[173][1]=16'hfff9,loc[173][2]=16'hfffd,loc[173][3]=16'h0000,loc[173][4]=16'h0008,loc[173][5]=16'hfff9,loc[173][6]=16'h0000,loc[173][7]=16'h0004,loc[173][8]=16'h0002,loc[173][9]=16'h000a,loc[173][10]=16'hfff9,loc[174][1]=16'h0001,loc[174][2]=16'h0000,loc[174][3]=16'h0008,loc[174][4]=16'hfffe,loc[174][5]=16'hfffe,loc[174][6]=16'h000a,loc[174][7]=16'hfff8,loc[174][8]=16'h0002,loc[174][9]=16'h0001,loc[174][10]=16'hfff8,loc[175][1]=16'h0000,loc[175][2]=16'h0002,loc[175][3]=16'h0004,loc[175][4]=16'hfffb,loc[175][5]=16'h0005,loc[175][6]=16'h0004,loc[175][7]=16'hfffb,loc[175][8]=16'h0005,loc[175][9]=16'hfff8,loc[175][10]=16'h0001,loc[176][1]=16'hfff6,loc[176][2]=16'hfffc,loc[176][3]=16'h0001,loc[176][4]=16'hfffa,loc[176][5]=16'h0003,loc[176][6]=16'hfff9,loc[176][7]=16'h0002,loc[176][8]=16'h0003,loc[176][9]=16'h000e,loc[176][10]=16'h000a,loc[177][1]=16'h000b,loc[177][2]=16'h000e,loc[177][3]=16'h000e,loc[177][4]=16'hfff7,loc[177][5]=16'h0005,loc[177][6]=16'hfff7,loc[177][7]=16'hfff4,loc[177][8]=16'hfffd,loc[177][9]=16'h0004,loc[177][10]=16'h0002,loc[178][1]=16'h0002,loc[178][2]=16'h0001,loc[178][3]=16'hfffb,loc[178][4]=16'hfff7,loc[178][5]=16'h0003,loc[178][6]=16'h0002,loc[178][7]=16'hfffb,loc[178][8]=16'h0019,loc[178][9]=16'hfff5,loc[178][10]=16'hfffe,loc[179][1]=16'h0005,loc[179][2]=16'hffff,loc[179][3]=16'hffff,loc[179][4]=16'hfffb,loc[179][5]=16'h0004,loc[179][6]=16'h000a,loc[179][7]=16'hfffe,loc[179][8]=16'hfffd,loc[179][9]=16'hfffe,loc[179][10]=16'hfffe,loc[180][1]=16'hfffe,loc[180][2]=16'hffff,loc[180][3]=16'h0001,loc[180][4]=16'hfffc,loc[180][5]=16'h0016,loc[180][6]=16'h0001,loc[180][7]=16'hfff3,loc[180][8]=16'hfff8,loc[180][9]=16'h0009,loc[180][10]=16'hffff,loc[181][1]=16'hfff8,loc[181][2]=16'h0000,loc[181][3]=16'h0002,loc[181][4]=16'hfffc,loc[181][5]=16'h0006,loc[181][6]=16'h0009,loc[181][7]=16'hfff4,loc[181][8]=16'hfffd,loc[181][9]=16'h0014,loc[181][10]=16'hfffa,loc[182][1]=16'h0002,loc[182][2]=16'hfffa,loc[182][3]=16'h0001,loc[182][4]=16'h0001,loc[182][5]=16'hfffd,loc[182][6]=16'hfffc,loc[182][7]=16'h0006,loc[182][8]=16'h000b,loc[182][9]=16'hffff,loc[182][10]=16'hfff9,loc[183][1]=16'h0006,loc[183][2]=16'h0002,loc[183][3]=16'h0002,loc[183][4]=16'hfffe,loc[183][5]=16'hfffd,loc[183][6]=16'h000b,loc[183][7]=16'hfffc,loc[183][8]=16'h0000,loc[183][9]=16'hfffe,loc[183][10]=16'hfffa,loc[184][1]=16'hfff9,loc[184][2]=16'h000e,loc[184][3]=16'hfffc,loc[184][4]=16'hfffd,loc[184][5]=16'hfff8,loc[184][6]=16'hfff4,loc[184][7]=16'h000e,loc[184][8]=16'h0005,loc[184][9]=16'h0006,loc[184][10]=16'h0001,loc[185][1]=16'hfffb,loc[185][2]=16'hfff6,loc[185][3]=16'h0004,loc[185][4]=16'hfff8,loc[185][5]=16'h0009,loc[185][6]=16'h0008,loc[185][7]=16'hffff,loc[185][8]=16'h0001,loc[185][9]=16'h0001,loc[185][10]=16'h0000,loc[186][1]=16'hffff,loc[186][2]=16'h0003,loc[186][3]=16'h000c,loc[186][4]=16'h0023,loc[186][5]=16'hfffb,loc[186][6]=16'hfffa,loc[186][7]=16'h0017,loc[186][8]=16'hfffb,loc[186][9]=16'hffda,loc[186][10]=16'hfff5,loc[187][1]=16'h0003,loc[187][2]=16'hffff,loc[187][3]=16'hfff7,loc[187][4]=16'hffff,loc[187][5]=16'hfffd,loc[187][6]=16'h0013,loc[187][7]=16'hfff8,loc[187][8]=16'h000e,loc[187][9]=16'hfff6,loc[187][10]=16'h0000,loc[188][1]=16'h001f,loc[188][2]=16'h0005,loc[188][3]=16'hfffa,loc[188][4]=16'hfffc,loc[188][5]=16'hfffe,loc[188][6]=16'h0000,loc[188][7]=16'hfff1,loc[188][8]=16'h0009,loc[188][9]=16'h0004,loc[188][10]=16'hfff0,loc[189][1]=16'hffff,loc[189][2]=16'h0002,loc[189][3]=16'h0008,loc[189][4]=16'h0005,loc[189][5]=16'h0001,loc[189][6]=16'hfff7,loc[189][7]=16'h0003,loc[189][8]=16'hfff8,loc[189][9]=16'hfff4,loc[189][10]=16'h000b,loc[190][1]=16'hfffe,loc[190][2]=16'hfff2,loc[190][3]=16'h0011,loc[190][4]=16'hfff9,loc[190][5]=16'h0003,loc[190][6]=16'hffeb,loc[190][7]=16'h0002,loc[190][8]=16'h0004,loc[190][9]=16'h0006,loc[190][10]=16'h0011,loc[191][1]=16'h0005,loc[191][2]=16'h0003,loc[191][3]=16'hfffd,loc[191][4]=16'h0005,loc[191][5]=16'h000b,loc[191][6]=16'h0004,loc[191][7]=16'hfff0,loc[191][8]=16'hfff8,loc[191][9]=16'h0006,loc[191][10]=16'hfffa,loc[192][1]=16'h0001,loc[192][2]=16'h0004,loc[192][3]=16'hfffc,loc[192][4]=16'h0005,loc[192][5]=16'hfffe,loc[192][6]=16'h0004,loc[192][7]=16'hfff9,loc[192][8]=16'hfffe,loc[192][9]=16'h000b,loc[192][10]=16'hfff7,loc[193][1]=16'h0001,loc[193][2]=16'h0015,loc[193][3]=16'hfff9,loc[193][4]=16'h0002,loc[193][5]=16'h0004,loc[193][6]=16'h0004,loc[193][7]=16'hffff,loc[193][8]=16'hffef,loc[193][9]=16'hfffc,loc[193][10]=16'h0003,loc[194][1]=16'hfffd,loc[194][2]=16'hfffa,loc[194][3]=16'h0003,loc[194][4]=16'h0002,loc[194][5]=16'h0002,loc[194][6]=16'hfffa,loc[194][7]=16'h0007,loc[194][8]=16'h0002,loc[194][9]=16'hfffe,loc[194][10]=16'h0002,loc[195][1]=16'hfff2,loc[195][2]=16'h0012,loc[195][3]=16'h0004,loc[195][4]=16'hfff6,loc[195][5]=16'h0021,loc[195][6]=16'hfff9,loc[195][7]=16'hfff9,loc[195][8]=16'hfff2,loc[195][9]=16'h0009,loc[195][10]=16'hfffc,loc[196][1]=16'hffff,loc[196][2]=16'h0002,loc[196][3]=16'hfffe,loc[196][4]=16'h0002,loc[196][5]=16'hfffe,loc[196][6]=16'h000e,loc[196][7]=16'hffff,loc[196][8]=16'h0003,loc[196][9]=16'hfff9,loc[196][10]=16'hfffc,loc[197][1]=16'h0004,loc[197][2]=16'h0001,loc[197][3]=16'hfffc,loc[197][4]=16'hfffd,loc[197][5]=16'h0005,loc[197][6]=16'h0004,loc[197][7]=16'h0003,loc[197][8]=16'hfffa,loc[197][9]=16'hffff,loc[197][10]=16'hfffc,loc[198][1]=16'h0008,loc[198][2]=16'hfff6,loc[198][3]=16'h0003,loc[198][4]=16'h0003,loc[198][5]=16'h0005,loc[198][6]=16'hffff,loc[198][7]=16'hfff8,loc[198][8]=16'h0003,loc[198][9]=16'h0001,loc[198][10]=16'hfffe,loc[199][1]=16'hffff,loc[199][2]=16'hfff6,loc[199][3]=16'h0002,loc[199][4]=16'hfffe,loc[199][5]=16'h0005,loc[199][6]=16'h0004,loc[199][7]=16'hfffb,loc[199][8]=16'h0004,loc[199][9]=16'h0003,loc[199][10]=16'hfffe,loc[200][1]=16'h0000,loc[200][2]=16'hfffa,loc[200][3]=16'h0002,loc[200][4]=16'hffff,loc[200][5]=16'h000a,loc[200][6]=16'hffff,loc[200][7]=16'h0003,loc[200][8]=16'hffff,loc[200][9]=16'h0002,loc[200][10]=16'hfffa,loc[201][1]=16'hfffe,loc[201][2]=16'hfff5,loc[201][3]=16'h0000,loc[201][4]=16'h0004,loc[201][5]=16'h0015,loc[201][6]=16'h0000,loc[201][7]=16'hfffd,loc[201][8]=16'hfff8,loc[201][9]=16'h0000,loc[201][10]=16'hffff,loc[202][1]=16'hfffa,loc[202][2]=16'hfff7,loc[202][3]=16'h0003,loc[202][4]=16'hffe6,loc[202][5]=16'hfff4,loc[202][6]=16'h0005,loc[202][7]=16'hfffc,loc[202][8]=16'h000e,loc[202][9]=16'h0009,loc[202][10]=16'h001c,loc[203][1]=16'h0005,loc[203][2]=16'h0008,loc[203][3]=16'hfffe,loc[203][4]=16'h0007,loc[203][5]=16'hfffb,loc[203][6]=16'hffff,loc[203][7]=16'h0007,loc[203][8]=16'h000c,loc[203][9]=16'hfffe,loc[203][10]=16'hffe5,loc[204][1]=16'hfffb,loc[204][2]=16'h0003,loc[204][3]=16'h0002,loc[204][4]=16'hfffa,loc[204][5]=16'hfffe,loc[204][6]=16'h0001,loc[204][7]=16'h0003,loc[204][8]=16'hffff,loc[204][9]=16'h0005,loc[204][10]=16'h0002,loc[205][1]=16'h0002,loc[205][2]=16'hfff7,loc[205][3]=16'h0007,loc[205][4]=16'h0000,loc[205][5]=16'h0004,loc[205][6]=16'h000c,loc[205][7]=16'h0001,loc[205][8]=16'h0004,loc[205][9]=16'hfff5,loc[205][10]=16'hfff8,loc[206][1]=16'hfffc,loc[206][2]=16'h0001,loc[206][3]=16'h0004,loc[206][4]=16'h0001,loc[206][5]=16'h0005,loc[206][6]=16'hfff8,loc[206][7]=16'h0006,loc[206][8]=16'hfff6,loc[206][9]=16'h0001,loc[206][10]=16'h0004,loc[207][1]=16'hfffb,loc[207][2]=16'hfff8,loc[207][3]=16'hfff7,loc[207][4]=16'h000e,loc[207][5]=16'h0004,loc[207][6]=16'h0005,loc[207][7]=16'h0002,loc[207][8]=16'hfffe,loc[207][9]=16'h0004,loc[207][10]=16'h0001,loc[208][1]=16'hfffa,loc[208][2]=16'h0000,loc[208][3]=16'hfffa,loc[208][4]=16'hfffb,loc[208][5]=16'h0002,loc[208][6]=16'h0002,loc[208][7]=16'h0001,loc[208][8]=16'h0003,loc[208][9]=16'h0006,loc[208][10]=16'h0007,loc[209][1]=16'hfffe,loc[209][2]=16'h0002,loc[209][3]=16'hfffc,loc[209][4]=16'h0005,loc[209][5]=16'h0003,loc[209][6]=16'hfff8,loc[209][7]=16'h0002,loc[209][8]=16'hfff2,loc[209][9]=16'h0009,loc[209][10]=16'h0003,loc[210][1]=16'h0004,loc[210][2]=16'hffff,loc[210][3]=16'h0004,loc[210][4]=16'h0001,loc[210][5]=16'h0001,loc[210][6]=16'hffff,loc[210][7]=16'h0003,loc[210][8]=16'hffff,loc[210][9]=16'hfff2,loc[210][10]=16'h0003,loc[211][1]=16'hffff,loc[211][2]=16'hfffa,loc[211][3]=16'hfffc,loc[211][4]=16'hffff,loc[211][5]=16'hfffa,loc[211][6]=16'hfffe,loc[211][7]=16'h0005,loc[211][8]=16'h000b,loc[211][9]=16'h0008,loc[211][10]=16'hfffd,loc[212][1]=16'hfff3,loc[212][2]=16'h0007,loc[212][3]=16'h000e,loc[212][4]=16'h0001,loc[212][5]=16'hfffe,loc[212][6]=16'hffff,loc[212][7]=16'h0005,loc[212][8]=16'h0002,loc[212][9]=16'hffea,loc[212][10]=16'h0005,loc[213][1]=16'h0000,loc[213][2]=16'h0006,loc[213][3]=16'h0001,loc[213][4]=16'hffff,loc[213][5]=16'h0004,loc[213][6]=16'h0000,loc[213][7]=16'hfff9,loc[213][8]=16'hfffa,loc[213][9]=16'h0005,loc[213][10]=16'h0003,loc[214][1]=16'hfffe,loc[214][2]=16'hfffb,loc[214][3]=16'h0006,loc[214][4]=16'h0005,loc[214][5]=16'hffff,loc[214][6]=16'h0004,loc[214][7]=16'hfffc,loc[214][8]=16'hfff9,loc[214][9]=16'h0002,loc[214][10]=16'h0003,loc[215][1]=16'hfffd,loc[215][2]=16'h0006,loc[215][3]=16'hfffb,loc[215][4]=16'h0006,loc[215][5]=16'hfffd,loc[215][6]=16'hffff,loc[215][7]=16'h0005,loc[215][8]=16'hfffb,loc[215][9]=16'hfffc,loc[215][10]=16'h0003,loc[216][1]=16'hfffa,loc[216][2]=16'hfffc,loc[216][3]=16'h0011,loc[216][4]=16'h000e,loc[216][5]=16'h0007,loc[216][6]=16'hfffa,loc[216][7]=16'h0007,loc[216][8]=16'hfff3,loc[216][9]=16'hfff9,loc[216][10]=16'hfff8,loc[217][1]=16'h0006,loc[217][2]=16'h0006,loc[217][3]=16'hfffa,loc[217][4]=16'h000e,loc[217][5]=16'h0000,loc[217][6]=16'hffff,loc[217][7]=16'h0000,loc[217][8]=16'hfffb,loc[217][9]=16'hfffc,loc[217][10]=16'hfffb,loc[218][1]=16'hffee,loc[218][2]=16'h0005,loc[218][3]=16'hfffc,loc[218][4]=16'hfffd,loc[218][5]=16'h0005,loc[218][6]=16'hfffe,loc[218][7]=16'h000d,loc[218][8]=16'h0003,loc[218][9]=16'hfff2,loc[218][10]=16'h0011,loc[219][1]=16'h0003,loc[219][2]=16'h0002,loc[219][3]=16'h0001,loc[219][4]=16'h0001,loc[219][5]=16'h0001,loc[219][6]=16'h000a,loc[219][7]=16'hfffd,loc[219][8]=16'hfffb,loc[219][9]=16'hfffd,loc[219][10]=16'hfffc,loc[220][1]=16'h0000,loc[220][2]=16'h0004,loc[220][3]=16'hfff5,loc[220][4]=16'hfffe,loc[220][5]=16'h0001,loc[220][6]=16'h0002,loc[220][7]=16'h0003,loc[220][8]=16'h0008,loc[220][9]=16'hfff9,loc[220][10]=16'h0001,loc[221][1]=16'h0001,loc[221][2]=16'hffed,loc[221][3]=16'h0005,loc[221][4]=16'h0003,loc[221][5]=16'h000b,loc[221][6]=16'hfffa,loc[221][7]=16'h0007,loc[221][8]=16'hffff,loc[221][9]=16'hfff4,loc[221][10]=16'h0007,loc[222][1]=16'hffff,loc[222][2]=16'h0001,loc[222][3]=16'hfff4,loc[222][4]=16'hffff,loc[222][5]=16'h0006,loc[222][6]=16'h0004,loc[222][7]=16'h0008,loc[222][8]=16'hfffa,loc[222][9]=16'hfffc,loc[222][10]=16'h0004,loc[223][1]=16'h0002,loc[223][2]=16'hfff5,loc[223][3]=16'hfffe,loc[223][4]=16'h0001,loc[223][5]=16'hfffc,loc[223][6]=16'hfff8,loc[223][7]=16'hfff2,loc[223][8]=16'h0014,loc[223][9]=16'h0011,loc[223][10]=16'h0002,loc[224][1]=16'hffff,loc[224][2]=16'hfffb,loc[224][3]=16'h000a,loc[224][4]=16'h0000,loc[224][5]=16'hffff,loc[224][6]=16'h0002,loc[224][7]=16'hffff,loc[224][8]=16'h0000,loc[224][9]=16'h0001,loc[224][10]=16'hffff,loc[225][1]=16'h0005,loc[225][2]=16'hffff,loc[225][3]=16'h0015,loc[225][4]=16'h0000,loc[225][5]=16'h0007,loc[225][6]=16'hffff,loc[225][7]=16'h0004,loc[225][8]=16'hfff7,loc[225][9]=16'hfff0,loc[225][10]=16'hfffb,loc[226][1]=16'h0005,loc[226][2]=16'h0001,loc[226][3]=16'hffff,loc[226][4]=16'h0004,loc[226][5]=16'h0008,loc[226][6]=16'h0000,loc[226][7]=16'hfff2,loc[226][8]=16'h0000,loc[226][9]=16'h0007,loc[226][10]=16'hfff6,loc[227][1]=16'hfff8,loc[227][2]=16'h0002,loc[227][3]=16'h0008,loc[227][4]=16'h0004,loc[227][5]=16'h0008,loc[227][6]=16'hfffe,loc[227][7]=16'hfff6,loc[227][8]=16'hffff,loc[227][9]=16'h0003,loc[227][10]=16'hffff,loc[228][1]=16'hfffa,loc[228][2]=16'h0001,loc[228][3]=16'hfffb,loc[228][4]=16'hffff,loc[228][5]=16'h0008,loc[228][6]=16'h0001,loc[228][7]=16'h0004,loc[228][8]=16'h0000,loc[228][9]=16'h0006,loc[228][10]=16'hfffa,loc[229][1]=16'hfffe,loc[229][2]=16'hfff6,loc[229][3]=16'h0001,loc[229][4]=16'h000a,loc[229][5]=16'h0011,loc[229][6]=16'hfffe,loc[229][7]=16'hffff,loc[229][8]=16'hfff6,loc[229][9]=16'h0006,loc[229][10]=16'hfffb,loc[230][1]=16'hfffd,loc[230][2]=16'h0004,loc[230][3]=16'hfffe,loc[230][4]=16'hfffc,loc[230][5]=16'h0003,loc[230][6]=16'h0000,loc[230][7]=16'h0005,loc[230][8]=16'hfffe,loc[230][9]=16'hfff4,loc[230][10]=16'h000b,loc[231][1]=16'hfffe,loc[231][2]=16'h0001,loc[231][3]=16'hfffe,loc[231][4]=16'hfffa,loc[231][5]=16'h0008,loc[231][6]=16'h0000,loc[231][7]=16'hfffe,loc[231][8]=16'hfffe,loc[231][9]=16'h0009,loc[231][10]=16'hfffd,loc[232][1]=16'hffff,loc[232][2]=16'hfff6,loc[232][3]=16'h0003,loc[232][4]=16'h0004,loc[232][5]=16'h000c,loc[232][6]=16'h0000,loc[232][7]=16'hffff,loc[232][8]=16'hfff7,loc[232][9]=16'hfff7,loc[232][10]=16'h000e,loc[233][1]=16'h0003,loc[233][2]=16'h0004,loc[233][3]=16'h0002,loc[233][4]=16'h000a,loc[233][5]=16'hfffb,loc[233][6]=16'h0007,loc[233][7]=16'hfff9,loc[233][8]=16'hfff7,loc[233][9]=16'hfff8,loc[233][10]=16'h0007,loc[234][1]=16'hfffe,loc[234][2]=16'hfffb,loc[234][3]=16'hfffa,loc[234][4]=16'hfffb,loc[234][5]=16'h0008,loc[234][6]=16'h0007,loc[234][7]=16'h0000,loc[234][8]=16'h0005,loc[234][9]=16'hffff,loc[234][10]=16'hfffe,loc[235][1]=16'h0001,loc[235][2]=16'h0001,loc[235][3]=16'hfffd,loc[235][4]=16'hfff5,loc[235][5]=16'hfff3,loc[235][6]=16'h0007,loc[235][7]=16'hfffe,loc[235][8]=16'h000c,loc[235][9]=16'hfffd,loc[235][10]=16'h000f,loc[236][1]=16'hfffe,loc[236][2]=16'h000e,loc[236][3]=16'hfffc,loc[236][4]=16'h0000,loc[236][5]=16'hfffe,loc[236][6]=16'h000c,loc[236][7]=16'hfffc,loc[236][8]=16'hfffa,loc[236][9]=16'hffff,loc[236][10]=16'hfffc,loc[237][1]=16'hfffe,loc[237][2]=16'hfffb,loc[237][3]=16'hfffe,loc[237][4]=16'h0002,loc[237][5]=16'hfffb,loc[237][6]=16'hfff7,loc[237][7]=16'h0005,loc[237][8]=16'h0001,loc[237][9]=16'h000f,loc[237][10]=16'hffff,loc[238][1]=16'h0003,loc[238][2]=16'h0003,loc[238][3]=16'hfffe,loc[238][4]=16'hfffb,loc[238][5]=16'h0001,loc[238][6]=16'h0006,loc[238][7]=16'hfffe,loc[238][8]=16'h0006,loc[238][9]=16'h0005,loc[238][10]=16'hfff8,loc[239][1]=16'hfffc,loc[239][2]=16'h0001,loc[239][3]=16'h0008,loc[239][4]=16'h0002,loc[239][5]=16'h0000,loc[239][6]=16'hfff9,loc[239][7]=16'h0002,loc[239][8]=16'h0002,loc[239][9]=16'h0000,loc[239][10]=16'hffff,loc[240][1]=16'hffff,loc[240][2]=16'h000a,loc[240][3]=16'h000d,loc[240][4]=16'hfffb,loc[240][5]=16'h0000,loc[240][6]=16'h0006,loc[240][7]=16'hfff0,loc[240][8]=16'hfffb,loc[240][9]=16'h0005,loc[240][10]=16'hfffe,loc[241][1]=16'h0001,loc[241][2]=16'h0009,loc[241][3]=16'h0006,loc[241][4]=16'h0001,loc[241][5]=16'hfffc,loc[241][6]=16'h0000,loc[241][7]=16'h0002,loc[241][8]=16'hfff3,loc[241][9]=16'hffee,loc[241][10]=16'h0012,loc[242][1]=16'hfffb,loc[242][2]=16'hffff,loc[242][3]=16'h0001,loc[242][4]=16'hfffc,loc[242][5]=16'h0004,loc[242][6]=16'h0004,loc[242][7]=16'hfffb,loc[242][8]=16'h0002,loc[242][9]=16'h0003,loc[242][10]=16'h0002,loc[243][1]=16'h001a,loc[243][2]=16'hfffe,loc[243][3]=16'hffec,loc[243][4]=16'hffe6,loc[243][5]=16'hfffa,loc[243][6]=16'hfff8,loc[243][7]=16'hffe8,loc[243][8]=16'h0018,loc[243][9]=16'h0002,loc[243][10]=16'h0021,loc[244][1]=16'h0000,loc[244][2]=16'h0013,loc[244][3]=16'hffff,loc[244][4]=16'h0001,loc[244][5]=16'h0005,loc[244][6]=16'hfff8,loc[244][7]=16'hfffe,loc[244][8]=16'hffee,loc[244][9]=16'h0001,loc[244][10]=16'h0007,loc[245][1]=16'hffff,loc[245][2]=16'hfff4,loc[245][3]=16'h0009,loc[245][4]=16'h0004,loc[245][5]=16'h0007,loc[245][6]=16'hfffd,loc[245][7]=16'h0001,loc[245][8]=16'hffff,loc[245][9]=16'h0005,loc[245][10]=16'hfffe,loc[246][1]=16'h0002,loc[246][2]=16'hfffd,loc[246][3]=16'hffff,loc[246][4]=16'h0004,loc[246][5]=16'h0005,loc[246][6]=16'h0004,loc[246][7]=16'h0004,loc[246][8]=16'hfffa,loc[246][9]=16'hfff9,loc[246][10]=16'h0003,loc[247][1]=16'hfffc,loc[247][2]=16'hfffb,loc[247][3]=16'hfffc,loc[247][4]=16'h0003,loc[247][5]=16'h0001,loc[247][6]=16'hfffc,loc[247][7]=16'h000d,loc[247][8]=16'hffff,loc[247][9]=16'h0004,loc[247][10]=16'hffff,loc[248][1]=16'hffff,loc[248][2]=16'hfffa,loc[248][3]=16'hfffd,loc[248][4]=16'h0000,loc[248][5]=16'hfffb,loc[248][6]=16'h0001,loc[248][7]=16'h0003,loc[248][8]=16'h0000,loc[248][9]=16'h0009,loc[248][10]=16'h0002,loc[249][1]=16'hfffd,loc[249][2]=16'h000e,loc[249][3]=16'hfff6,loc[249][4]=16'hfffd,loc[249][5]=16'h0000,loc[249][6]=16'h0006,loc[249][7]=16'hfffe,loc[249][8]=16'hfffc,loc[249][9]=16'h0009,loc[249][10]=16'hfffe,loc[250][1]=16'hfffa,loc[250][2]=16'hfffe,loc[250][3]=16'hfffe,loc[250][4]=16'hffff,loc[250][5]=16'h0006,loc[250][6]=16'h000a,loc[250][7]=16'hfff8,loc[250][8]=16'h0001,loc[250][9]=16'h0009,loc[250][10]=16'hfffa,loc[251][1]=16'h0006,loc[251][2]=16'h0006,loc[251][3]=16'hfffd,loc[251][4]=16'h0000,loc[251][5]=16'hfff9,loc[251][6]=16'hffea,loc[251][7]=16'h0005,loc[251][8]=16'h0010,loc[251][9]=16'hffea,loc[251][10]=16'h0014,loc[252][1]=16'h0004,loc[252][2]=16'h0015,loc[252][3]=16'h0001,loc[252][4]=16'h0000,loc[252][5]=16'hfff6,loc[252][6]=16'hfff3,loc[252][7]=16'h000a,loc[252][8]=16'h0002,loc[252][9]=16'hfff8,loc[252][10]=16'hfffe,loc[253][1]=16'hffee,loc[253][2]=16'hfffd,loc[253][3]=16'h0003,loc[253][4]=16'hffed,loc[253][5]=16'hfffa,loc[253][6]=16'h0015,loc[253][7]=16'hffec,loc[253][8]=16'h000b,loc[253][9]=16'h0015,loc[253][10]=16'h000c,loc[254][1]=16'h0006,loc[254][2]=16'h0009,loc[254][3]=16'hfff3,loc[254][4]=16'h0001,loc[254][5]=16'hfff8,loc[254][6]=16'h0000,loc[254][7]=16'h0004,loc[254][8]=16'h0004,loc[254][9]=16'h0003,loc[254][10]=16'hffff,loc[255][1]=16'hffff,loc[255][2]=16'h0000,loc[255][3]=16'hfff8,loc[255][4]=16'h0004,loc[255][5]=16'hfffb,loc[255][6]=16'h0003,loc[255][7]=16'h0001,loc[255][8]=16'hffff,loc[255][9]=16'h0007,loc[255][10]=16'h0002,loc[256][1]=16'h0005,loc[256][2]=16'h0001,loc[256][3]=16'h0003,loc[256][4]=16'h0001,loc[256][5]=16'h0007,loc[256][6]=16'h0008,loc[256][7]=16'hfffb,loc[256][8]=16'h0005,loc[256][9]=16'hffea,loc[256][10]=16'hffff,loc[257][1]=16'h0000,loc[257][2]=16'h0000,loc[257][3]=16'h0000,loc[257][4]=16'h0000,loc[257][5]=16'h0000,loc[257][6]=16'h0000,loc[257][7]=16'h0000,loc[257][8]=16'h0000,loc[257][9]=16'h0000,loc[257][10]=16'h0000,loc[258][1]=16'h0009,loc[258][2]=16'h0008,loc[258][3]=16'h0007,loc[258][4]=16'hfffd,loc[258][5]=16'hffff,loc[258][6]=16'hfffc,loc[258][7]=16'h0000,loc[258][8]=16'h0001,loc[258][9]=16'hffed,loc[258][10]=16'h0003,loc[259][1]=16'hffff,loc[259][2]=16'h0001,loc[259][3]=16'h0000,loc[259][4]=16'h0004,loc[259][5]=16'h0002,loc[259][6]=16'h0000,loc[259][7]=16'hfffc,loc[259][8]=16'h0003,loc[259][9]=16'hfffc,loc[259][10]=16'h0004,loc[260][1]=16'hfffa,loc[260][2]=16'h000a,loc[260][3]=16'h0000,loc[260][4]=16'h0006,loc[260][5]=16'hfffb,loc[260][6]=16'hfffd,loc[260][7]=16'h000c,loc[260][8]=16'hffff,loc[260][9]=16'hfff9,loc[260][10]=16'hffff,loc[261][1]=16'h0009,loc[261][2]=16'hffff,loc[261][3]=16'h000b,loc[261][4]=16'hfff5,loc[261][5]=16'h0003,loc[261][6]=16'h0002,loc[261][7]=16'hfffc,loc[261][8]=16'h0001,loc[261][9]=16'hfffb,loc[261][10]=16'hfffb,loc[262][1]=16'h0002,loc[262][2]=16'h0004,loc[262][3]=16'h0004,loc[262][4]=16'hfffd,loc[262][5]=16'hfffe,loc[262][6]=16'hfffe,loc[262][7]=16'hfffb,loc[262][8]=16'h0002,loc[262][9]=16'h0005,loc[262][10]=16'hfffb,loc[263][1]=16'hffff,loc[263][2]=16'hfff9,loc[263][3]=16'h000a,loc[263][4]=16'h0003,loc[263][5]=16'hfffc,loc[263][6]=16'hfffb,loc[263][7]=16'hfffd,loc[263][8]=16'h0000,loc[263][9]=16'h0002,loc[263][10]=16'h0006,loc[264][1]=16'hfffd,loc[264][2]=16'h0002,loc[264][3]=16'hfff0,loc[264][4]=16'h0004,loc[264][5]=16'h000d,loc[264][6]=16'hfffc,loc[264][7]=16'hfffa,loc[264][8]=16'hfffc,loc[264][9]=16'h0017,loc[264][10]=16'hfff6,loc[265][1]=16'hfff9,loc[265][2]=16'h000f,loc[265][3]=16'h0010,loc[265][4]=16'hfffd,loc[265][5]=16'h0001,loc[265][6]=16'h0004,loc[265][7]=16'hfff5,loc[265][8]=16'hfff9,loc[265][9]=16'hfff6,loc[265][10]=16'h0004,loc[266][1]=16'hfffe,loc[266][2]=16'h0000,loc[266][3]=16'h0003,loc[266][4]=16'h0000,loc[266][5]=16'h0000,loc[266][6]=16'h0002,loc[266][7]=16'h0001,loc[266][8]=16'hfff3,loc[266][9]=16'h000e,loc[266][10]=16'hfffd,loc[267][1]=16'hfffb,loc[267][2]=16'h0004,loc[267][3]=16'h0004,loc[267][4]=16'h0007,loc[267][5]=16'hfffe,loc[267][6]=16'hfff8,loc[267][7]=16'h0006,loc[267][8]=16'h0001,loc[267][9]=16'hfff9,loc[267][10]=16'hfffd,loc[268][1]=16'hfffc,loc[268][2]=16'h0008,loc[268][3]=16'hfffd,loc[268][4]=16'hfffd,loc[268][5]=16'h0003,loc[268][6]=16'hfffc,loc[268][7]=16'h0000,loc[268][8]=16'hfffd,loc[268][9]=16'h0002,loc[268][10]=16'h0005,loc[269][1]=16'h0004,loc[269][2]=16'hffff,loc[269][3]=16'h0007,loc[269][4]=16'h0000,loc[269][5]=16'h0003,loc[269][6]=16'h0001,loc[269][7]=16'hfffb,loc[269][8]=16'hffff,loc[269][9]=16'h0001,loc[269][10]=16'hfff9,loc[270][1]=16'h0000,loc[270][2]=16'h0000,loc[270][3]=16'hffff,loc[270][4]=16'hfffb,loc[270][5]=16'h0006,loc[270][6]=16'hffff,loc[270][7]=16'hfffb,loc[270][8]=16'h0006,loc[270][9]=16'h0000,loc[270][10]=16'h0004,loc[271][1]=16'h0005,loc[271][2]=16'hffff,loc[271][3]=16'h0001,loc[271][4]=16'h0009,loc[271][5]=16'hfffb,loc[271][6]=16'hfff9,loc[271][7]=16'h0004,loc[271][8]=16'hfffd,loc[271][9]=16'hfffd,loc[271][10]=16'h0002,loc[272][1]=16'h0001,loc[272][2]=16'hffff,loc[272][3]=16'h0009,loc[272][4]=16'h0004,loc[272][5]=16'h0005,loc[272][6]=16'h0001,loc[272][7]=16'hffff,loc[272][8]=16'hfffc,loc[272][9]=16'hfffd,loc[272][10]=16'hfffb,loc[273][1]=16'h0000,loc[273][2]=16'h0005,loc[273][3]=16'hfff8,loc[273][4]=16'hfffd,loc[273][5]=16'hfffd,loc[273][6]=16'h000c,loc[273][7]=16'hfffe,loc[273][8]=16'h0006,loc[273][9]=16'h0007,loc[273][10]=16'hfff0,loc[274][1]=16'h0005,loc[274][2]=16'h0004,loc[274][3]=16'hfff6,loc[274][4]=16'h0008,loc[274][5]=16'hfffc,loc[274][6]=16'hfffd,loc[274][7]=16'h0000,loc[274][8]=16'h0002,loc[274][9]=16'hfff7,loc[274][10]=16'h0005,loc[275][1]=16'hfff5,loc[275][2]=16'hfff7,loc[275][3]=16'h000a,loc[275][4]=16'h0006,loc[275][5]=16'h0002,loc[275][6]=16'hfffd,loc[275][7]=16'h0008,loc[275][8]=16'hfffc,loc[275][9]=16'hfff6,loc[275][10]=16'h000a,loc[276][1]=16'h0008,loc[276][2]=16'h0012,loc[276][3]=16'h0009,loc[276][4]=16'hfffd,loc[276][5]=16'hfff5,loc[276][6]=16'hffff,loc[276][7]=16'hfff7,loc[276][8]=16'hfff6,loc[276][9]=16'hfff5,loc[276][10]=16'h0012,loc[277][1]=16'hfff5,loc[277][2]=16'h0003,loc[277][3]=16'h0000,loc[277][4]=16'h0006,loc[277][5]=16'h0004,loc[277][6]=16'hfff9,loc[277][7]=16'h0003,loc[277][8]=16'h0003,loc[277][9]=16'hffff,loc[277][10]=16'h0004,loc[278][1]=16'h0008,loc[278][2]=16'hfffb,loc[278][3]=16'h0007,loc[278][4]=16'hfff2,loc[278][5]=16'h0000,loc[278][6]=16'h0000,loc[278][7]=16'hfffd,loc[278][8]=16'h000d,loc[278][9]=16'h0000,loc[278][10]=16'hffff,loc[279][1]=16'h0003,loc[279][2]=16'h0001,loc[279][3]=16'h0006,loc[279][4]=16'hfffd,loc[279][5]=16'hfffd,loc[279][6]=16'h0002,loc[279][7]=16'hfff0,loc[279][8]=16'hfffd,loc[279][9]=16'h0009,loc[279][10]=16'h0003,loc[280][1]=16'hffff,loc[280][2]=16'hfffb,loc[280][3]=16'h0009,loc[280][4]=16'h0005,loc[280][5]=16'hffff,loc[280][6]=16'h0000,loc[280][7]=16'h0008,loc[280][8]=16'hfffa,loc[280][9]=16'h0002,loc[280][10]=16'hfffd,loc[281][1]=16'hfffd,loc[281][2]=16'hfff5,loc[281][3]=16'hfffc,loc[281][4]=16'h0002,loc[281][5]=16'h0003,loc[281][6]=16'h0001,loc[281][7]=16'hfffc,loc[281][8]=16'h000d,loc[281][9]=16'hfffe,loc[281][10]=16'h0007,loc[282][1]=16'h0001,loc[282][2]=16'h0007,loc[282][3]=16'h0009,loc[282][4]=16'hfffe,loc[282][5]=16'h0008,loc[282][6]=16'hffff,loc[282][7]=16'hfffc,loc[282][8]=16'hfffa,loc[282][9]=16'hfffd,loc[282][10]=16'hfffc,loc[283][1]=16'hfffb,loc[283][2]=16'hffed,loc[283][3]=16'h000b,loc[283][4]=16'hfff2,loc[283][5]=16'h0000,loc[283][6]=16'h0003,loc[283][7]=16'h0004,loc[283][8]=16'h0013,loc[283][9]=16'h0003,loc[283][10]=16'hfffb,loc[284][1]=16'hfffc,loc[284][2]=16'hfffd,loc[284][3]=16'h0007,loc[284][4]=16'h0000,loc[284][5]=16'hfffc,loc[284][6]=16'hfff9,loc[284][7]=16'h0006,loc[284][8]=16'h0006,loc[284][9]=16'hfff1,loc[284][10]=16'h000f,loc[285][1]=16'hfff1,loc[285][2]=16'h0006,loc[285][3]=16'hfff6,loc[285][4]=16'hffe6,loc[285][5]=16'h000f,loc[285][6]=16'h0017,loc[285][7]=16'h000d,loc[285][8]=16'hffe4,loc[285][9]=16'h0013,loc[285][10]=16'h000c,loc[286][1]=16'h0001,loc[286][2]=16'h0000,loc[286][3]=16'hffff,loc[286][4]=16'h0004,loc[286][5]=16'h0000,loc[286][6]=16'hffff,loc[286][7]=16'h0001,loc[286][8]=16'h0001,loc[286][9]=16'hfff7,loc[286][10]=16'h0006,loc[287][1]=16'hfffa,loc[287][2]=16'hfff9,loc[287][3]=16'h0004,loc[287][4]=16'h0000,loc[287][5]=16'h000c,loc[287][6]=16'hfff6,loc[287][7]=16'h0004,loc[287][8]=16'h0001,loc[287][9]=16'hfffc,loc[287][10]=16'h0009,loc[288][1]=16'hfffc,loc[288][2]=16'hfffe,loc[288][3]=16'hfffe,loc[288][4]=16'hfffb,loc[288][5]=16'h0002,loc[288][6]=16'hfffe,loc[288][7]=16'h0001,loc[288][8]=16'h0008,loc[288][9]=16'h0004,loc[288][10]=16'h0001,loc[289][1]=16'h0000,loc[289][2]=16'h0000,loc[289][3]=16'hfff9,loc[289][4]=16'h000b,loc[289][5]=16'hfff6,loc[289][6]=16'h0014,loc[289][7]=16'hfffd,loc[289][8]=16'hfff0,loc[289][9]=16'h0006,loc[289][10]=16'h0004,loc[290][1]=16'hfff4,loc[290][2]=16'hfffa,loc[290][3]=16'h0006,loc[290][4]=16'h0006,loc[290][5]=16'h000b,loc[290][6]=16'hfff6,loc[290][7]=16'hfffc,loc[290][8]=16'h0011,loc[290][9]=16'hfffd,loc[290][10]=16'hfffd,loc[291][1]=16'h000b,loc[291][2]=16'hfff0,loc[291][3]=16'h0003,loc[291][4]=16'hfffd,loc[291][5]=16'hfffc,loc[291][6]=16'hfffd,loc[291][7]=16'h000d,loc[291][8]=16'h0001,loc[291][9]=16'h0008,loc[291][10]=16'hfff3,loc[292][1]=16'hfffb,loc[292][2]=16'h0001,loc[292][3]=16'hfffe,loc[292][4]=16'hfffd,loc[292][5]=16'hfff8,loc[292][6]=16'hfff6,loc[292][7]=16'h000d,loc[292][8]=16'h0000,loc[292][9]=16'hffff,loc[292][10]=16'h000e,loc[293][1]=16'hfffb,loc[293][2]=16'h0002,loc[293][3]=16'h0001,loc[293][4]=16'hfffe,loc[293][5]=16'hfffb,loc[293][6]=16'hfffd,loc[293][7]=16'h000b,loc[293][8]=16'h0002,loc[293][9]=16'hfff3,loc[293][10]=16'h000d,loc[294][1]=16'h0004,loc[294][2]=16'hfffd,loc[294][3]=16'h0006,loc[294][4]=16'h0007,loc[294][5]=16'hfff7,loc[294][6]=16'hfff9,loc[294][7]=16'h0002,loc[294][8]=16'h0007,loc[294][9]=16'hfffd,loc[294][10]=16'hfff9,loc[295][1]=16'hfff5,loc[295][2]=16'h0007,loc[295][3]=16'h0011,loc[295][4]=16'hfffd,loc[295][5]=16'hfff3,loc[295][6]=16'h0023,loc[295][7]=16'hfffa,loc[295][8]=16'h0003,loc[295][9]=16'h0002,loc[295][10]=16'hffeb,loc[296][1]=16'hfffc,loc[296][2]=16'hffff,loc[296][3]=16'hfff4,loc[296][4]=16'h000a,loc[296][5]=16'hfffe,loc[296][6]=16'hfff2,loc[296][7]=16'h000a,loc[296][8]=16'hfffa,loc[296][9]=16'h0011,loc[296][10]=16'h0002,loc[297][1]=16'hfffc,loc[297][2]=16'hfffc,loc[297][3]=16'h0000,loc[297][4]=16'h0002,loc[297][5]=16'h0001,loc[297][6]=16'hfff5,loc[297][7]=16'h0006,loc[297][8]=16'hfffd,loc[297][9]=16'h000d,loc[297][10]=16'hffff,loc[298][1]=16'h0001,loc[298][2]=16'h000a,loc[298][3]=16'hfffd,loc[298][4]=16'hfffb,loc[298][5]=16'hfffc,loc[298][6]=16'h0004,loc[298][7]=16'h0001,loc[298][8]=16'h0004,loc[298][9]=16'hfffe,loc[298][10]=16'h0002,loc[299][1]=16'hfffb,loc[299][2]=16'h0005,loc[299][3]=16'hfffb,loc[299][4]=16'hfffc,loc[299][5]=16'hfffc,loc[299][6]=16'hfffa,loc[299][7]=16'hffff,loc[299][8]=16'h0005,loc[299][9]=16'h000c,loc[299][10]=16'h0000,loc[300][1]=16'h0000,loc[300][2]=16'h000a,loc[300][3]=16'h0002,loc[300][4]=16'h0001,loc[300][5]=16'hfff3,loc[300][6]=16'hfff4,loc[300][7]=16'h0005,loc[300][8]=16'h0005,loc[300][9]=16'h000e,loc[300][10]=16'hfff2,loc[301][1]=16'h0002,loc[301][2]=16'h0012,loc[301][3]=16'hfff4,loc[301][4]=16'h000c,loc[301][5]=16'hfffc,loc[301][6]=16'h0008,loc[301][7]=16'h0004,loc[301][8]=16'hffef,loc[301][9]=16'h0001,loc[301][10]=16'hfff6,loc[302][1]=16'hfffc,loc[302][2]=16'hfff4,loc[302][3]=16'hfffd,loc[302][4]=16'hfff5,loc[302][5]=16'h000a,loc[302][6]=16'hfffb,loc[302][7]=16'hfffc,loc[302][8]=16'h0010,loc[302][9]=16'h0004,loc[302][10]=16'h000f,loc[303][1]=16'hfffb,loc[303][2]=16'h000e,loc[303][3]=16'hfffd,loc[303][4]=16'h000c,loc[303][5]=16'hfffc,loc[303][6]=16'h0001,loc[303][7]=16'hffff,loc[303][8]=16'hfff1,loc[303][9]=16'hfffd,loc[303][10]=16'hffff,loc[304][1]=16'h0003,loc[304][2]=16'h000a,loc[304][3]=16'h0005,loc[304][4]=16'hfff7,loc[304][5]=16'h0005,loc[304][6]=16'h0009,loc[304][7]=16'hfffd,loc[304][8]=16'hfff5,loc[304][9]=16'hfff8,loc[304][10]=16'h0003,loc[305][1]=16'h0007,loc[305][2]=16'h0008,loc[305][3]=16'h0000,loc[305][4]=16'hfffa,loc[305][5]=16'hffd8,loc[305][6]=16'hfff9,loc[305][7]=16'h0006,loc[305][8]=16'h000d,loc[305][9]=16'h0004,loc[305][10]=16'h000c,loc[306][1]=16'hfff8,loc[306][2]=16'h0001,loc[306][3]=16'h0006,loc[306][4]=16'h0012,loc[306][5]=16'hfffa,loc[306][6]=16'hfffc,loc[306][7]=16'h0008,loc[306][8]=16'hfffd,loc[306][9]=16'hfff3,loc[306][10]=16'h0005,loc[307][1]=16'h0007,loc[307][2]=16'hfffe,loc[307][3]=16'hfffc,loc[307][4]=16'h0004,loc[307][5]=16'hfff5,loc[307][6]=16'hfffd,loc[307][7]=16'h0003,loc[307][8]=16'h000b,loc[307][9]=16'h0000,loc[307][10]=16'h0006,loc[308][1]=16'h0000,loc[308][2]=16'h0000,loc[308][3]=16'h0000,loc[308][4]=16'h0000,loc[308][5]=16'h0000,loc[308][6]=16'h0000,loc[308][7]=16'h0000,loc[308][8]=16'h0000,loc[308][9]=16'h0000,loc[308][10]=16'h0000,loc[309][1]=16'hfffe,loc[309][2]=16'h0002,loc[309][3]=16'hfffc,loc[309][4]=16'hfff5,loc[309][5]=16'hfffa,loc[309][6]=16'h0003,loc[309][7]=16'h0002,loc[309][8]=16'h000b,loc[309][9]=16'h0005,loc[309][10]=16'h0004,loc[310][1]=16'hfff8,loc[310][2]=16'hfff8,loc[310][3]=16'hfff6,loc[310][4]=16'hfff8,loc[310][5]=16'h0007,loc[310][6]=16'hffff,loc[310][7]=16'h0009,loc[310][8]=16'h0001,loc[310][9]=16'hfffc,loc[310][10]=16'h0014,loc[311][1]=16'hfffb,loc[311][2]=16'h0007,loc[311][3]=16'hfffd,loc[311][4]=16'h0006,loc[311][5]=16'hfffd,loc[311][6]=16'hfff8,loc[311][7]=16'h0013,loc[311][8]=16'hfffb,loc[311][9]=16'hfffa,loc[311][10]=16'hfffc,loc[312][1]=16'hfffe,loc[312][2]=16'h0003,loc[312][3]=16'hfffb,loc[312][4]=16'h0003,loc[312][5]=16'h0004,loc[312][6]=16'hfff6,loc[312][7]=16'hfffc,loc[312][8]=16'h0004,loc[312][9]=16'h0005,loc[312][10]=16'h0001,loc[313][1]=16'hfffd,loc[313][2]=16'h0008,loc[313][3]=16'hfffa,loc[313][4]=16'hfff5,loc[313][5]=16'h0002,loc[313][6]=16'h001b,loc[313][7]=16'hfffe,loc[313][8]=16'hfff2,loc[313][9]=16'h0009,loc[313][10]=16'h0000,loc[314][1]=16'h0005,loc[314][2]=16'h0004,loc[314][3]=16'h0005,loc[314][4]=16'hfffd,loc[314][5]=16'hfffc,loc[314][6]=16'h000d,loc[314][7]=16'hfffb,loc[314][8]=16'hffff,loc[314][9]=16'hfffd,loc[314][10]=16'hfff4,loc[315][1]=16'hfffb,loc[315][2]=16'h0000,loc[315][3]=16'h0008,loc[315][4]=16'h0000,loc[315][5]=16'h0006,loc[315][6]=16'h0008,loc[315][7]=16'hffff,loc[315][8]=16'h0003,loc[315][9]=16'hfff6,loc[315][10]=16'hfff9,loc[316][1]=16'h0002,loc[316][2]=16'hfff8,loc[316][3]=16'h0004,loc[316][4]=16'hfffc,loc[316][5]=16'hfffd,loc[316][6]=16'hffff,loc[316][7]=16'h0004,loc[316][8]=16'h0002,loc[316][9]=16'hfffe,loc[316][10]=16'h0005,loc[317][1]=16'hfffe,loc[317][2]=16'hfffd,loc[317][3]=16'h000b,loc[317][4]=16'h0006,loc[317][5]=16'hfff9,loc[317][6]=16'hfffd,loc[317][7]=16'h000c,loc[317][8]=16'hfffc,loc[317][9]=16'hfff9,loc[317][10]=16'h0000,loc[318][1]=16'hfffe,loc[318][2]=16'hfffd,loc[318][3]=16'h000c,loc[318][4]=16'hfffc,loc[318][5]=16'h0005,loc[318][6]=16'hfffb,loc[318][7]=16'h0001,loc[318][8]=16'hfff2,loc[318][9]=16'hffff,loc[318][10]=16'h0009,loc[319][1]=16'h0002,loc[319][2]=16'hfff4,loc[319][3]=16'h0001,loc[319][4]=16'h0009,loc[319][5]=16'h0004,loc[319][6]=16'h0003,loc[319][7]=16'hffff,loc[319][8]=16'hfffc,loc[319][9]=16'h0006,loc[319][10]=16'hfff8,loc[320][1]=16'hffff,loc[320][2]=16'h0002,loc[320][3]=16'hfff5,loc[320][4]=16'hfffb,loc[320][5]=16'h000f,loc[320][6]=16'hfffe,loc[320][7]=16'hfffc,loc[320][8]=16'h0001,loc[320][9]=16'hfff5,loc[320][10]=16'h0010,loc[321][1]=16'hffff,loc[321][2]=16'hfffa,loc[321][3]=16'h0006,loc[321][4]=16'hfffc,loc[321][5]=16'hfffd,loc[321][6]=16'h000c,loc[321][7]=16'hfffa,loc[321][8]=16'h0006,loc[321][9]=16'hfffd,loc[321][10]=16'hffff,loc[322][1]=16'hfffb,loc[322][2]=16'hfff4,loc[322][3]=16'h0009,loc[322][4]=16'hfffc,loc[322][5]=16'hffff,loc[322][6]=16'h0002,loc[322][7]=16'h0002,loc[322][8]=16'h0002,loc[322][9]=16'hffff,loc[322][10]=16'h0007,loc[323][1]=16'hfffa,loc[323][2]=16'hfff8,loc[323][3]=16'h0008,loc[323][4]=16'hffff,loc[323][5]=16'h0006,loc[323][6]=16'hfffd,loc[323][7]=16'h0000,loc[323][8]=16'h000f,loc[323][9]=16'h0001,loc[323][10]=16'hfff7,loc[324][1]=16'h0002,loc[324][2]=16'hfffe,loc[324][3]=16'hfff9,loc[324][4]=16'hfff6,loc[324][5]=16'hfffd,loc[324][6]=16'h0004,loc[324][7]=16'h0003,loc[324][8]=16'h0001,loc[324][9]=16'h0001,loc[324][10]=16'h0008,loc[325][1]=16'hffff,loc[325][2]=16'h0000,loc[325][3]=16'h0009,loc[325][4]=16'hfff7,loc[325][5]=16'h0004,loc[325][6]=16'h0010,loc[325][7]=16'hfff9,loc[325][8]=16'h0001,loc[325][9]=16'hfffc,loc[325][10]=16'hfffc,loc[326][1]=16'hfff9,loc[326][2]=16'hfffd,loc[326][3]=16'hfff1,loc[326][4]=16'h0009,loc[326][5]=16'h0008,loc[326][6]=16'h0000,loc[326][7]=16'h0005,loc[326][8]=16'h0005,loc[326][9]=16'hfffa,loc[326][10]=16'h0006,loc[327][1]=16'hffff,loc[327][2]=16'h0003,loc[327][3]=16'hfffc,loc[327][4]=16'hffff,loc[327][5]=16'h0000,loc[327][6]=16'h0006,loc[327][7]=16'h0000,loc[327][8]=16'hffff,loc[327][9]=16'h0006,loc[327][10]=16'hfff9,loc[328][1]=16'h0002,loc[328][2]=16'hfff9,loc[328][3]=16'h0000,loc[328][4]=16'h0005,loc[328][5]=16'hfffd,loc[328][6]=16'hfff7,loc[328][7]=16'h0009,loc[328][8]=16'hffff,loc[328][9]=16'h0001,loc[328][10]=16'hfffd,loc[329][1]=16'hfffa,loc[329][2]=16'h0008,loc[329][3]=16'hfffb,loc[329][4]=16'h0002,loc[329][5]=16'h0002,loc[329][6]=16'h0008,loc[329][7]=16'h0002,loc[329][8]=16'hfff5,loc[329][9]=16'h0001,loc[329][10]=16'h0000,loc[330][1]=16'hffff,loc[330][2]=16'hfffe,loc[330][3]=16'h0002,loc[330][4]=16'hfff6,loc[330][5]=16'h0001,loc[330][6]=16'hfffe,loc[330][7]=16'hfff7,loc[330][8]=16'h000f,loc[330][9]=16'h0004,loc[330][10]=16'h0001,loc[331][1]=16'h0002,loc[331][2]=16'hfff5,loc[331][3]=16'h0005,loc[331][4]=16'hfffd,loc[331][5]=16'h0006,loc[331][6]=16'h0003,loc[331][7]=16'h0005,loc[331][8]=16'h0001,loc[331][9]=16'hfffe,loc[331][10]=16'hfffc,loc[332][1]=16'h0001,loc[332][2]=16'h0001,loc[332][3]=16'hfffb,loc[332][4]=16'h0005,loc[332][5]=16'h0000,loc[332][6]=16'hfffb,loc[332][7]=16'h0002,loc[332][8]=16'hfffe,loc[332][9]=16'h0005,loc[332][10]=16'h0002,loc[333][1]=16'h0000,loc[333][2]=16'hffff,loc[333][3]=16'h0003,loc[333][4]=16'h0003,loc[333][5]=16'h0002,loc[333][6]=16'h0003,loc[333][7]=16'h0000,loc[333][8]=16'hfffa,loc[333][9]=16'hfff8,loc[333][10]=16'h0001,loc[334][1]=16'hffec,loc[334][2]=16'h0000,loc[334][3]=16'hffeb,loc[334][4]=16'h0017,loc[334][5]=16'hfff7,loc[334][6]=16'h0008,loc[334][7]=16'hfffd,loc[334][8]=16'hfff6,loc[334][9]=16'h0015,loc[334][10]=16'h0002,loc[335][1]=16'h0005,loc[335][2]=16'h000c,loc[335][3]=16'h0003,loc[335][4]=16'hfff2,loc[335][5]=16'hfffe,loc[335][6]=16'h0002,loc[335][7]=16'h0000,loc[335][8]=16'hfff6,loc[335][9]=16'h0008,loc[335][10]=16'hfffc,loc[336][1]=16'h0004,loc[336][2]=16'hfff7,loc[336][3]=16'h0004,loc[336][4]=16'hffff,loc[336][5]=16'h0003,loc[336][6]=16'hfff5,loc[336][7]=16'h0002,loc[336][8]=16'h0006,loc[336][9]=16'hfffc,loc[336][10]=16'h0004,loc[337][1]=16'h0001,loc[337][2]=16'h0003,loc[337][3]=16'hfff9,loc[337][4]=16'h0006,loc[337][5]=16'hfffc,loc[337][6]=16'hfffd,loc[337][7]=16'h0001,loc[337][8]=16'h0000,loc[337][9]=16'h0005,loc[337][10]=16'h0002,loc[338][1]=16'h0000,loc[338][2]=16'h0016,loc[338][3]=16'hfffc,loc[338][4]=16'hfff3,loc[338][5]=16'hfffe,loc[338][6]=16'h0001,loc[338][7]=16'h0005,loc[338][8]=16'hfffc,loc[338][9]=16'hfffe,loc[338][10]=16'hffff,loc[339][1]=16'h0000,loc[339][2]=16'hfffb,loc[339][3]=16'h0003,loc[339][4]=16'hfff8,loc[339][5]=16'hfff9,loc[339][6]=16'h0005,loc[339][7]=16'hfffc,loc[339][8]=16'h0007,loc[339][9]=16'h0006,loc[339][10]=16'h0001,loc[340][1]=16'hffff,loc[340][2]=16'h0003,loc[340][3]=16'hfff6,loc[340][4]=16'hffff,loc[340][5]=16'h0006,loc[340][6]=16'h000d,loc[340][7]=16'hfffc,loc[340][8]=16'h0003,loc[340][9]=16'hfff4,loc[340][10]=16'h0008,loc[341][1]=16'hfffe,loc[341][2]=16'hfffb,loc[341][3]=16'hfffc,loc[341][4]=16'h0002,loc[341][5]=16'h0004,loc[341][6]=16'h0001,loc[341][7]=16'h0000,loc[341][8]=16'h0001,loc[341][9]=16'h0005,loc[341][10]=16'h0001,loc[342][1]=16'h0003,loc[342][2]=16'h000f,loc[342][3]=16'h0006,loc[342][4]=16'hffff,loc[342][5]=16'hfff6,loc[342][6]=16'h0004,loc[342][7]=16'hfff8,loc[342][8]=16'h0003,loc[342][9]=16'hfffc,loc[342][10]=16'hfffb,loc[343][1]=16'h0003,loc[343][2]=16'h0001,loc[343][3]=16'hfffe,loc[343][4]=16'hfff9,loc[343][5]=16'hfffb,loc[343][6]=16'hfff3,loc[343][7]=16'h0000,loc[343][8]=16'h0007,loc[343][9]=16'h0002,loc[343][10]=16'h000c,loc[344][1]=16'hfffb,loc[344][2]=16'h000b,loc[344][3]=16'h0000,loc[344][4]=16'hfff5,loc[344][5]=16'h0001,loc[344][6]=16'h0007,loc[344][7]=16'hffff,loc[344][8]=16'h0003,loc[344][9]=16'hfff7,loc[344][10]=16'h0007,loc[345][1]=16'hfff9,loc[345][2]=16'hfffe,loc[345][3]=16'h000c,loc[345][4]=16'h0011,loc[345][5]=16'hfff6,loc[345][6]=16'h0007,loc[345][7]=16'h0004,loc[345][8]=16'hfffa,loc[345][9]=16'hfff3,loc[345][10]=16'h0002,loc[346][1]=16'h0004,loc[346][2]=16'h0006,loc[346][3]=16'h0004,loc[346][4]=16'hfffe,loc[346][5]=16'hfffa,loc[346][6]=16'hfffd,loc[346][7]=16'hfffd,loc[346][8]=16'hfffe,loc[346][9]=16'h000b,loc[346][10]=16'hfff6,loc[347][1]=16'hfffd,loc[347][2]=16'h0004,loc[347][3]=16'hfffe,loc[347][4]=16'h0002,loc[347][5]=16'hfffc,loc[347][6]=16'hfffc,loc[347][7]=16'hfffd,loc[347][8]=16'h0002,loc[347][9]=16'h000a,loc[347][10]=16'hfffd,loc[348][1]=16'h0004,loc[348][2]=16'h0002,loc[348][3]=16'h0007,loc[348][4]=16'h0003,loc[348][5]=16'h0001,loc[348][6]=16'hfffd,loc[348][7]=16'hfffc,loc[348][8]=16'hfffc,loc[348][9]=16'h0000,loc[348][10]=16'hfffa,loc[349][1]=16'hfffa,loc[349][2]=16'hffff,loc[349][3]=16'h0003,loc[349][4]=16'h0000,loc[349][5]=16'hfffd,loc[349][6]=16'hfffd,loc[349][7]=16'h0003,loc[349][8]=16'hfffe,loc[349][9]=16'h0005,loc[349][10]=16'h0000,loc[350][1]=16'hfffe,loc[350][2]=16'h0009,loc[350][3]=16'hfffe,loc[350][4]=16'hfffc,loc[350][5]=16'h0009,loc[350][6]=16'h000b,loc[350][7]=16'hfff4,loc[350][8]=16'hfff9,loc[350][9]=16'hfffd,loc[350][10]=16'h0002,loc[351][1]=16'h000c,loc[351][2]=16'h0020,loc[351][3]=16'h000a,loc[351][4]=16'hfff4,loc[351][5]=16'hfff7,loc[351][6]=16'hfffd,loc[351][7]=16'h0009,loc[351][8]=16'h0001,loc[351][9]=16'hffea,loc[351][10]=16'hfff9,loc[352][1]=16'h0004,loc[352][2]=16'h0008,loc[352][3]=16'h0007,loc[352][4]=16'hfff9,loc[352][5]=16'hfff9,loc[352][6]=16'h0001,loc[352][7]=16'hfffe,loc[352][8]=16'hfffd,loc[352][9]=16'h0002,loc[352][10]=16'hfffe,loc[353][1]=16'hffff,loc[353][2]=16'hfff7,loc[353][3]=16'hfffc,loc[353][4]=16'hfffe,loc[353][5]=16'h0001,loc[353][6]=16'hffff,loc[353][7]=16'hffff,loc[353][8]=16'h0006,loc[353][9]=16'h000a,loc[353][10]=16'h0004,loc[354][1]=16'h0000,loc[354][2]=16'h0003,loc[354][3]=16'h0003,loc[354][4]=16'h0001,loc[354][5]=16'hfffd,loc[354][6]=16'h0002,loc[354][7]=16'hfff3,loc[354][8]=16'h0001,loc[354][9]=16'h0009,loc[354][10]=16'hfffc,loc[355][1]=16'hfffc,loc[355][2]=16'h0005,loc[355][3]=16'h0008,loc[355][4]=16'hfff6,loc[355][5]=16'h000c,loc[355][6]=16'h0009,loc[355][7]=16'hfff1,loc[355][8]=16'h0009,loc[355][9]=16'h0004,loc[355][10]=16'hfff1,loc[356][1]=16'h0006,loc[356][2]=16'hfffc,loc[356][3]=16'hfffd,loc[356][4]=16'hfffd,loc[356][5]=16'hfffd,loc[356][6]=16'hfff7,loc[356][7]=16'h0002,loc[356][8]=16'h000a,loc[356][9]=16'h0003,loc[356][10]=16'h0002,loc[357][1]=16'h0001,loc[357][2]=16'hfffd,loc[357][3]=16'h0006,loc[357][4]=16'h0007,loc[357][5]=16'h0003,loc[357][6]=16'hfff6,loc[357][7]=16'hfff8,loc[357][8]=16'h0000,loc[357][9]=16'h0003,loc[357][10]=16'h0000,loc[358][1]=16'h0005,loc[358][2]=16'h0007,loc[358][3]=16'h0000,loc[358][4]=16'hffff,loc[358][5]=16'h0000,loc[358][6]=16'h0006,loc[358][7]=16'hfff5,loc[358][8]=16'hfffa,loc[358][9]=16'h0006,loc[358][10]=16'hfffd,loc[359][1]=16'hfff5,loc[359][2]=16'hffe9,loc[359][3]=16'h000e,loc[359][4]=16'h0008,loc[359][5]=16'h0010,loc[359][6]=16'hfff2,loc[359][7]=16'h0002,loc[359][8]=16'h000f,loc[359][9]=16'hfffd,loc[359][10]=16'hfffe,loc[360][1]=16'hfffc,loc[360][2]=16'hfff8,loc[360][3]=16'hfffc,loc[360][4]=16'hfffe,loc[360][5]=16'h0004,loc[360][6]=16'h0007,loc[360][7]=16'h0000,loc[360][8]=16'h0004,loc[360][9]=16'hfffb,loc[360][10]=16'h000c,loc[361][1]=16'hfff2,loc[361][2]=16'hfff8,loc[361][3]=16'hfffa,loc[361][4]=16'hffe8,loc[361][5]=16'h0001,loc[361][6]=16'h0007,loc[361][7]=16'h0005,loc[361][8]=16'h0012,loc[361][9]=16'h000b,loc[361][10]=16'h0012,loc[362][1]=16'hfffe,loc[362][2]=16'h0004,loc[362][3]=16'hfff3,loc[362][4]=16'hfff9,loc[362][5]=16'hfffa,loc[362][6]=16'h000b,loc[362][7]=16'h000e,loc[362][8]=16'h0001,loc[362][9]=16'hfff8,loc[362][10]=16'h0007,loc[363][1]=16'hfffb,loc[363][2]=16'h0002,loc[363][3]=16'hfffd,loc[363][4]=16'h000c,loc[363][5]=16'h0001,loc[363][6]=16'hfff7,loc[363][7]=16'h0002,loc[363][8]=16'h0000,loc[363][9]=16'h0002,loc[363][10]=16'hfffe,loc[364][1]=16'h0003,loc[364][2]=16'hfff7,loc[364][3]=16'h0010,loc[364][4]=16'h0002,loc[364][5]=16'h0003,loc[364][6]=16'hfffb,loc[364][7]=16'hfff9,loc[364][8]=16'h0000,loc[364][9]=16'hfffb,loc[364][10]=16'hffff,loc[365][1]=16'h000b,loc[365][2]=16'hffff,loc[365][3]=16'h0001,loc[365][4]=16'h0000,loc[365][5]=16'hfffa,loc[365][6]=16'h000c,loc[365][7]=16'hfff8,loc[365][8]=16'hfff9,loc[365][9]=16'h0000,loc[365][10]=16'h0002,loc[366][1]=16'hfffc,loc[366][2]=16'hfffe,loc[366][3]=16'hfffe,loc[366][4]=16'h0014,loc[366][5]=16'h0006,loc[366][6]=16'h0003,loc[366][7]=16'h0005,loc[366][8]=16'hfff9,loc[366][9]=16'hfff2,loc[366][10]=16'hfffe,loc[367][1]=16'h0002,loc[367][2]=16'hfffd,loc[367][3]=16'h0003,loc[367][4]=16'h0005,loc[367][5]=16'hfffb,loc[367][6]=16'hfff9,loc[367][7]=16'h0001,loc[367][8]=16'hfff2,loc[367][9]=16'h0013,loc[367][10]=16'hffff,loc[368][1]=16'hfffb,loc[368][2]=16'h0005,loc[368][3]=16'h0007,loc[368][4]=16'hfff4,loc[368][5]=16'hffff,loc[368][6]=16'h000b,loc[368][7]=16'hfff6,loc[368][8]=16'h0007,loc[368][9]=16'h000b,loc[368][10]=16'hfff2,loc[369][1]=16'h0007,loc[369][2]=16'hfffc,loc[369][3]=16'hfffe,loc[369][4]=16'hfffa,loc[369][5]=16'hfffc,loc[369][6]=16'hffff,loc[369][7]=16'hfffa,loc[369][8]=16'hfffd,loc[369][9]=16'hfffe,loc[369][10]=16'h0012,loc[370][1]=16'h0006,loc[370][2]=16'h0000,loc[370][3]=16'h0001,loc[370][4]=16'h0003,loc[370][5]=16'h0007,loc[370][6]=16'h0006,loc[370][7]=16'h0000,loc[370][8]=16'hfffc,loc[370][9]=16'hfff3,loc[370][10]=16'hfffa,loc[371][1]=16'hfff9,loc[371][2]=16'hfffc,loc[371][3]=16'h0003,loc[371][4]=16'h0004,loc[371][5]=16'h0008,loc[371][6]=16'hfffb,loc[371][7]=16'hffff,loc[371][8]=16'hffff,loc[371][9]=16'h0000,loc[371][10]=16'h0002,loc[372][1]=16'hffff,loc[372][2]=16'hfffc,loc[372][3]=16'hffff,loc[372][4]=16'h0003,loc[372][5]=16'h0006,loc[372][6]=16'h0000,loc[372][7]=16'h0004,loc[372][8]=16'hfffc,loc[372][9]=16'hfffd,loc[372][10]=16'h0000,loc[373][1]=16'h0019,loc[373][2]=16'hffc6,loc[373][3]=16'hffc8,loc[373][4]=16'hffdc,loc[373][5]=16'h0017,loc[373][6]=16'h0078,loc[373][7]=16'hffde,loc[373][8]=16'h0075,loc[373][9]=16'hfff1,loc[373][10]=16'hffbd,loc[374][1]=16'h0003,loc[374][2]=16'h0004,loc[374][3]=16'hffff,loc[374][4]=16'hfffb,loc[374][5]=16'h0001,loc[374][6]=16'h0002,loc[374][7]=16'hfff7,loc[374][8]=16'h0005,loc[374][9]=16'h0003,loc[374][10]=16'hffff,loc[375][1]=16'hffff,loc[375][2]=16'hfff9,loc[375][3]=16'h0002,loc[375][4]=16'hffff,loc[375][5]=16'h0006,loc[375][6]=16'hfffa,loc[375][7]=16'h0003,loc[375][8]=16'h000c,loc[375][9]=16'hfffe,loc[375][10]=16'hffff,loc[376][1]=16'hfff5,loc[376][2]=16'h0003,loc[376][3]=16'hfffb,loc[376][4]=16'h0002,loc[376][5]=16'hffff,loc[376][6]=16'h0002,loc[376][7]=16'h0002,loc[376][8]=16'h0002,loc[376][9]=16'h0006,loc[376][10]=16'h0003,loc[377][1]=16'hfffb,loc[377][2]=16'h0006,loc[377][3]=16'h0000,loc[377][4]=16'h0001,loc[377][5]=16'hfff9,loc[377][6]=16'hfffe,loc[377][7]=16'h000b,loc[377][8]=16'hfffe,loc[377][9]=16'h0006,loc[377][10]=16'hfff8,loc[378][1]=16'hfff9,loc[378][2]=16'h0003,loc[378][3]=16'h0004,loc[378][4]=16'hfffb,loc[378][5]=16'hfffc,loc[378][6]=16'hfffc,loc[378][7]=16'h000b,loc[378][8]=16'hfff7,loc[378][9]=16'h0001,loc[378][10]=16'h0010,loc[379][1]=16'h0003,loc[379][2]=16'hfffe,loc[379][3]=16'h0002,loc[379][4]=16'hfffc,loc[379][5]=16'h0004,loc[379][6]=16'hfffe,loc[379][7]=16'hfffe,loc[379][8]=16'h0000,loc[379][9]=16'h0007,loc[379][10]=16'hfffd,loc[380][1]=16'h0002,loc[380][2]=16'hffff,loc[380][3]=16'h000d,loc[380][4]=16'h0006,loc[380][5]=16'h000b,loc[380][6]=16'h0001,loc[380][7]=16'h0000,loc[380][8]=16'hfff7,loc[380][9]=16'hfffa,loc[380][10]=16'hfff5,loc[381][1]=16'hfff5,loc[381][2]=16'hfffe,loc[381][3]=16'hfffb,loc[381][4]=16'h0003,loc[381][5]=16'h0001,loc[381][6]=16'h000e,loc[381][7]=16'h0000,loc[381][8]=16'h0005,loc[381][9]=16'h0002,loc[381][10]=16'hfffc,loc[382][1]=16'hfffe,loc[382][2]=16'h0004,loc[382][3]=16'h000b,loc[382][4]=16'hfff6,loc[382][5]=16'hfffd,loc[382][6]=16'h0000,loc[382][7]=16'h0002,loc[382][8]=16'h0003,loc[382][9]=16'hfff8,loc[382][10]=16'h0007,loc[383][1]=16'h0005,loc[383][2]=16'h0006,loc[383][3]=16'hfff2,loc[383][4]=16'h0016,loc[383][5]=16'hffff,loc[383][6]=16'h0000,loc[383][7]=16'hfffc,loc[383][8]=16'hfff7,loc[383][9]=16'h0005,loc[383][10]=16'hfffb,loc[384][1]=16'h0001,loc[384][2]=16'h002b,loc[384][3]=16'h0005,loc[384][4]=16'h0007,loc[384][5]=16'hfffc,loc[384][6]=16'hffff,loc[384][7]=16'h0013,loc[384][8]=16'hffd6,loc[384][9]=16'hffef,loc[384][10]=16'hfff4,loc[385][1]=16'h0004,loc[385][2]=16'hfffe,loc[385][3]=16'h0004,loc[385][4]=16'hffff,loc[385][5]=16'hfff9,loc[385][6]=16'h0000,loc[385][7]=16'hfffe,loc[385][8]=16'hffff,loc[385][9]=16'h0000,loc[385][10]=16'h0005,loc[386][1]=16'hfffd,loc[386][2]=16'hfffc,loc[386][3]=16'hfffa,loc[386][4]=16'h0001,loc[386][5]=16'h0007,loc[386][6]=16'h0012,loc[386][7]=16'hfffd,loc[386][8]=16'hfffe,loc[386][9]=16'h0000,loc[386][10]=16'hfff9,loc[387][1]=16'hffff,loc[387][2]=16'h0002,loc[387][3]=16'hfff9,loc[387][4]=16'hfff6,loc[387][5]=16'h0005,loc[387][6]=16'h0001,loc[387][7]=16'h0003,loc[387][8]=16'h0001,loc[387][9]=16'hfffd,loc[387][10]=16'h0009,loc[388][1]=16'hfffb,loc[388][2]=16'h0000,loc[388][3]=16'h0004,loc[388][4]=16'hffef,loc[388][5]=16'h0007,loc[388][6]=16'h0003,loc[388][7]=16'hffff,loc[388][8]=16'h0004,loc[388][9]=16'hffff,loc[388][10]=16'h0006,loc[389][1]=16'h0005,loc[389][2]=16'hfffd,loc[389][3]=16'hfffc,loc[389][4]=16'hfff8,loc[389][5]=16'hfffb,loc[389][6]=16'hfffc,loc[389][7]=16'h0004,loc[389][8]=16'h0009,loc[389][9]=16'h0000,loc[389][10]=16'h0001,loc[390][1]=16'hfffd,loc[390][2]=16'hfffd,loc[390][3]=16'h0004,loc[390][4]=16'h0004,loc[390][5]=16'h000a,loc[390][6]=16'h0005,loc[390][7]=16'hffff,loc[390][8]=16'hfff6,loc[390][9]=16'h0001,loc[390][10]=16'hfff9,loc[391][1]=16'h0000,loc[391][2]=16'hfffe,loc[391][3]=16'hfff6,loc[391][4]=16'h0008,loc[391][5]=16'h0000,loc[391][6]=16'h0003,loc[391][7]=16'h0000,loc[391][8]=16'hffff,loc[391][9]=16'h0005,loc[391][10]=16'hfffc,loc[392][1]=16'h0004,loc[392][2]=16'hfff4,loc[392][3]=16'hfffb,loc[392][4]=16'h0004,loc[392][5]=16'h0001,loc[392][6]=16'h0014,loc[392][7]=16'hfffb,loc[392][8]=16'h000a,loc[392][9]=16'hfffb,loc[392][10]=16'hfffb,loc[393][1]=16'h0001,loc[393][2]=16'h0005,loc[393][3]=16'h0001,loc[393][4]=16'hfffe,loc[393][5]=16'hfffa,loc[393][6]=16'hffff,loc[393][7]=16'h0008,loc[393][8]=16'hfffc,loc[393][9]=16'h0006,loc[393][10]=16'hfff7,loc[394][1]=16'h0004,loc[394][2]=16'h0000,loc[394][3]=16'hfffe,loc[394][4]=16'h0007,loc[394][5]=16'h0000,loc[394][6]=16'hfff9,loc[394][7]=16'h0003,loc[394][8]=16'hfff8,loc[394][9]=16'h0000,loc[394][10]=16'h0003,loc[395][1]=16'hfffd,loc[395][2]=16'hfffa,loc[395][3]=16'hfffe,loc[395][4]=16'hfffa,loc[395][5]=16'h0010,loc[395][6]=16'h0005,loc[395][7]=16'h0002,loc[395][8]=16'hffff,loc[395][9]=16'hfffa,loc[395][10]=16'h0002,loc[396][1]=16'hfffc,loc[396][2]=16'hfff8,loc[396][3]=16'hfffd,loc[396][4]=16'hfffc,loc[396][5]=16'h0005,loc[396][6]=16'h0003,loc[396][7]=16'hfffe,loc[396][8]=16'h0004,loc[396][9]=16'h0002,loc[396][10]=16'h0005,loc[397][1]=16'h0014,loc[397][2]=16'h0026,loc[397][3]=16'hffe6,loc[397][4]=16'hfff5,loc[397][5]=16'h0019,loc[397][6]=16'hffd9,loc[397][7]=16'h0001,loc[397][8]=16'hffd9,loc[397][9]=16'h0006,loc[397][10]=16'h0032,loc[398][1]=16'h0005,loc[398][2]=16'h000b,loc[398][3]=16'h0004,loc[398][4]=16'h0003,loc[398][5]=16'hfffc,loc[398][6]=16'h0009,loc[398][7]=16'h0008,loc[398][8]=16'hfff5,loc[398][9]=16'hfff1,loc[398][10]=16'hfff7,loc[399][1]=16'h0015,loc[399][2]=16'h0016,loc[399][3]=16'hffdd,loc[399][4]=16'hfffc,loc[399][5]=16'h0026,loc[399][6]=16'hffd4,loc[399][7]=16'hfff7,loc[399][8]=16'h0019,loc[399][9]=16'hffe0,loc[399][10]=16'h002b,loc[400][1]=16'hfff8,loc[400][2]=16'hfffa,loc[400][3]=16'hfffd,loc[400][4]=16'h0019,loc[400][5]=16'hfffd,loc[400][6]=16'hfffe,loc[400][7]=16'h0009,loc[400][8]=16'hfffd,loc[400][9]=16'hfffb,loc[400][10]=16'h0001,loc[401][1]=16'h0007,loc[401][2]=16'h0007,loc[401][3]=16'hffff,loc[401][4]=16'hfffb,loc[401][5]=16'hfffc,loc[401][6]=16'h0004,loc[401][7]=16'hfff8,loc[401][8]=16'h0003,loc[401][9]=16'hfffa,loc[401][10]=16'h0006,loc[402][1]=16'h0003,loc[402][2]=16'h0009,loc[402][3]=16'hfff5,loc[402][4]=16'h000b,loc[402][5]=16'hffff,loc[402][6]=16'hfff4,loc[402][7]=16'hfff5,loc[402][8]=16'hfffb,loc[402][9]=16'hffff,loc[402][10]=16'h0010,loc[403][1]=16'hfff4,loc[403][2]=16'hfff8,loc[403][3]=16'hfffd,loc[403][4]=16'h0009,loc[403][5]=16'hfffd,loc[403][6]=16'hfffc,loc[403][7]=16'h0009,loc[403][8]=16'h0006,loc[403][9]=16'h000b,loc[403][10]=16'hfff8,loc[404][1]=16'hfffe,loc[404][2]=16'hfff6,loc[404][3]=16'h0003,loc[404][4]=16'hffff,loc[404][5]=16'h0003,loc[404][6]=16'h0001,loc[404][7]=16'hffff,loc[404][8]=16'h000d,loc[404][9]=16'hfffd,loc[404][10]=16'hfffd,loc[405][1]=16'h0001,loc[405][2]=16'hfff9,loc[405][3]=16'h000b,loc[405][4]=16'hfffd,loc[405][5]=16'h0005,loc[405][6]=16'hfffe,loc[405][7]=16'hfffa,loc[405][8]=16'hfffa,loc[405][9]=16'h0014,loc[405][10]=16'hfff0,loc[406][1]=16'h0005,loc[406][2]=16'h0005,loc[406][3]=16'h0006,loc[406][4]=16'h000c,loc[406][5]=16'h0004,loc[406][6]=16'hfff9,loc[406][7]=16'hfffd,loc[406][8]=16'hffff,loc[406][9]=16'hfff1,loc[406][10]=16'hfffc,loc[407][1]=16'h0008,loc[407][2]=16'hfffb,loc[407][3]=16'hfffa,loc[407][4]=16'h0005,loc[407][5]=16'h0003,loc[407][6]=16'hfff5,loc[407][7]=16'hfff8,loc[407][8]=16'h000c,loc[407][9]=16'h0009,loc[407][10]=16'hfffc,loc[408][1]=16'hfff9,loc[408][2]=16'h0009,loc[408][3]=16'h000e,loc[408][4]=16'hfffa,loc[408][5]=16'h0006,loc[408][6]=16'hfffc,loc[408][7]=16'h0000,loc[408][8]=16'hfff6,loc[408][9]=16'hfff6,loc[408][10]=16'h0006,loc[409][1]=16'hffff,loc[409][2]=16'h0002,loc[409][3]=16'hfffd,loc[409][4]=16'h0001,loc[409][5]=16'h000d,loc[409][6]=16'h0006,loc[409][7]=16'hfff9,loc[409][8]=16'hfff7,loc[409][9]=16'h0009,loc[409][10]=16'hfff4,loc[410][1]=16'h0001,loc[410][2]=16'h0010,loc[410][3]=16'hfffe,loc[410][4]=16'hfffc,loc[410][5]=16'hfffb,loc[410][6]=16'h0006,loc[410][7]=16'hfff8,loc[410][8]=16'hfffb,loc[410][9]=16'h0002,loc[410][10]=16'h0001,loc[411][1]=16'h0002,loc[411][2]=16'h0000,loc[411][3]=16'hfff9,loc[411][4]=16'h0008,loc[411][5]=16'hfff1,loc[411][6]=16'hfff4,loc[411][7]=16'h0013,loc[411][8]=16'h0002,loc[411][9]=16'h0008,loc[411][10]=16'hfffb,loc[412][1]=16'hffff,loc[412][2]=16'hfffe,loc[412][3]=16'h0005,loc[412][4]=16'h0005,loc[412][5]=16'h0002,loc[412][6]=16'hfffe,loc[412][7]=16'hffff,loc[412][8]=16'hffff,loc[412][9]=16'hffff,loc[412][10]=16'hfffe,loc[413][1]=16'h0002,loc[413][2]=16'hfff2,loc[413][3]=16'h0006,loc[413][4]=16'h000e,loc[413][5]=16'h0000,loc[413][6]=16'h0002,loc[413][7]=16'h0001,loc[413][8]=16'h0001,loc[413][9]=16'hfffe,loc[413][10]=16'hfff5,loc[414][1]=16'h000a,loc[414][2]=16'hfffd,loc[414][3]=16'hffff,loc[414][4]=16'hfff9,loc[414][5]=16'hfffc,loc[414][6]=16'h0004,loc[414][7]=16'h0000,loc[414][8]=16'h0010,loc[414][9]=16'hfff5,loc[414][10]=16'hffff,loc[415][1]=16'h0002,loc[415][2]=16'hfffc,loc[415][3]=16'h000a,loc[415][4]=16'h0004,loc[415][5]=16'hffff,loc[415][6]=16'hfffa,loc[415][7]=16'hfff4,loc[415][8]=16'h000a,loc[415][9]=16'h0008,loc[415][10]=16'hfff7,loc[416][1]=16'h0004,loc[416][2]=16'h0008,loc[416][3]=16'h0001,loc[416][4]=16'hffed,loc[416][5]=16'hfffd,loc[416][6]=16'h000e,loc[416][7]=16'hfffa,loc[416][8]=16'h0009,loc[416][9]=16'hfffe,loc[416][10]=16'hfffc,loc[417][1]=16'hffe7,loc[417][2]=16'h0018,loc[417][3]=16'hfff2,loc[417][4]=16'h0005,loc[417][5]=16'hffef,loc[417][6]=16'h0017,loc[417][7]=16'h000b,loc[417][8]=16'hfff1,loc[417][9]=16'h000c,loc[417][10]=16'hfff0,loc[418][1]=16'h0002,loc[418][2]=16'hfffc,loc[418][3]=16'h0001,loc[418][4]=16'h0000,loc[418][5]=16'h0001,loc[418][6]=16'h0006,loc[418][7]=16'h0002,loc[418][8]=16'hffff,loc[418][9]=16'h0002,loc[418][10]=16'hfff7,loc[419][1]=16'hfff4,loc[419][2]=16'hfff2,loc[419][3]=16'hffff,loc[419][4]=16'h0002,loc[419][5]=16'hfff5,loc[419][6]=16'h0016,loc[419][7]=16'hfff7,loc[419][8]=16'h0023,loc[419][9]=16'h0004,loc[419][10]=16'hffef,loc[420][1]=16'hfffc,loc[420][2]=16'h0004,loc[420][3]=16'h0004,loc[420][4]=16'h0003,loc[420][5]=16'h0000,loc[420][6]=16'hfff5,loc[420][7]=16'h0003,loc[420][8]=16'hfffc,loc[420][9]=16'hfff8,loc[420][10]=16'h000a;

    always@(loc[1][1] or addr) begin
        case(addr)
            1:begin W21 = {loc[1][1],loc[1][2],loc[1][3],loc[1][4],loc[1][5],loc[1][6],loc[1][7],loc[1][8],loc[1][9],loc[1][10]};end	
            2:begin W21 = {loc[2][1],loc[2][2],loc[2][3],loc[2][4],loc[2][5],loc[2][6],loc[2][7],loc[2][8],loc[2][9],loc[2][10]};end
            3:begin W21 = {loc[3][1],loc[3][2],loc[3][3],loc[3][4],loc[3][5],loc[3][6],loc[3][7],loc[3][8],loc[3][9],loc[3][10]};end
            4:begin W21 = {loc[4][1],loc[4][2],loc[4][3],loc[4][4],loc[4][5],loc[4][6],loc[4][7],loc[4][8],loc[4][9],loc[4][10]};end
            5:begin W21 = {loc[5][1],loc[5][2],loc[5][3],loc[5][4],loc[5][5],loc[5][6],loc[5][7],loc[5][8],loc[5][9],loc[5][10]};end
            6:begin W21 = {loc[6][1],loc[6][2],loc[6][3],loc[6][4],loc[6][5],loc[6][6],loc[6][7],loc[6][8],loc[6][9],loc[6][10]};end
            7:begin W21 = {loc[7][1],loc[7][2],loc[7][3],loc[7][4],loc[7][5],loc[7][6],loc[7][7],loc[7][8],loc[7][9],loc[7][10]};end
            8:begin W21 = {loc[8][1],loc[8][2],loc[8][3],loc[8][4],loc[8][5],loc[8][6],loc[8][7],loc[8][8],loc[8][9],loc[8][10]};end
            9:begin W21 = {loc[9][1],loc[9][2],loc[9][3],loc[9][4],loc[9][5],loc[9][6],loc[9][7],loc[9][8],loc[9][9],loc[9][10]};end
            10:begin W21 = {loc[10][1],loc[10][2],loc[10][3],loc[10][4],loc[10][5],loc[10][6],loc[10][7],loc[10][8],loc[10][9],loc[10][10]};end
            11:begin W21 = {loc[11][1],loc[11][2],loc[11][3],loc[11][4],loc[11][5],loc[11][6],loc[11][7],loc[11][8],loc[11][9],loc[11][10]};end
            12:begin W21 = {loc[12][1],loc[12][2],loc[12][3],loc[12][4],loc[12][5],loc[12][6],loc[12][7],loc[12][8],loc[12][9],loc[12][10]};end
            13:begin W21 = {loc[13][1],loc[13][2],loc[13][3],loc[13][4],loc[13][5],loc[13][6],loc[13][7],loc[13][8],loc[13][9],loc[13][10]};end
            14:begin W21 = {loc[14][1],loc[14][2],loc[14][3],loc[14][4],loc[14][5],loc[14][6],loc[14][7],loc[14][8],loc[14][9],loc[14][10]};end
            15:begin W21 = {loc[15][1],loc[15][2],loc[15][3],loc[15][4],loc[15][5],loc[15][6],loc[15][7],loc[15][8],loc[15][9],loc[15][10]};end
            16:begin W21 = {loc[16][1],loc[16][2],loc[16][3],loc[16][4],loc[16][5],loc[16][6],loc[16][7],loc[16][8],loc[16][9],loc[16][10]};end
            17:begin W21 = {loc[17][1],loc[17][2],loc[17][3],loc[17][4],loc[17][5],loc[17][6],loc[17][7],loc[17][8],loc[17][9],loc[17][10]};end
            18:begin W21 = {loc[18][1],loc[18][2],loc[18][3],loc[18][4],loc[18][5],loc[18][6],loc[18][7],loc[18][8],loc[18][9],loc[18][10]};end
            19:begin W21 = {loc[19][1],loc[19][2],loc[19][3],loc[19][4],loc[19][5],loc[19][6],loc[19][7],loc[19][8],loc[19][9],loc[19][10]};end
            20:begin W21 = {loc[20][1],loc[20][2],loc[20][3],loc[20][4],loc[20][5],loc[20][6],loc[20][7],loc[20][8],loc[20][9],loc[20][10]};end
            21:begin W21 = {loc[21][1],loc[21][2],loc[21][3],loc[21][4],loc[21][5],loc[21][6],loc[21][7],loc[21][8],loc[21][9],loc[21][10]};end
            22:begin W21 = {loc[22][1],loc[22][2],loc[22][3],loc[22][4],loc[22][5],loc[22][6],loc[22][7],loc[22][8],loc[22][9],loc[22][10]};end
            23:begin W21 = {loc[23][1],loc[23][2],loc[23][3],loc[23][4],loc[23][5],loc[23][6],loc[23][7],loc[23][8],loc[23][9],loc[23][10]};end
            24:begin W21 = {loc[24][1],loc[24][2],loc[24][3],loc[24][4],loc[24][5],loc[24][6],loc[24][7],loc[24][8],loc[24][9],loc[24][10]};end
            25:begin W21 = {loc[25][1],loc[25][2],loc[25][3],loc[25][4],loc[25][5],loc[25][6],loc[25][7],loc[25][8],loc[25][9],loc[25][10]};end
            26:begin W21 = {loc[26][1],loc[26][2],loc[26][3],loc[26][4],loc[26][5],loc[26][6],loc[26][7],loc[26][8],loc[26][9],loc[26][10]};end
            27:begin W21 = {loc[27][1],loc[27][2],loc[27][3],loc[27][4],loc[27][5],loc[27][6],loc[27][7],loc[27][8],loc[27][9],loc[27][10]};end
            28:begin W21 = {loc[28][1],loc[28][2],loc[28][3],loc[28][4],loc[28][5],loc[28][6],loc[28][7],loc[28][8],loc[28][9],loc[28][10]};end
            29:begin W21 = {loc[29][1],loc[29][2],loc[29][3],loc[29][4],loc[29][5],loc[29][6],loc[29][7],loc[29][8],loc[29][9],loc[29][10]};end
            30:begin W21 = {loc[30][1],loc[30][2],loc[30][3],loc[30][4],loc[30][5],loc[30][6],loc[30][7],loc[30][8],loc[30][9],loc[30][10]};end
            31:begin W21 = {loc[31][1],loc[31][2],loc[31][3],loc[31][4],loc[31][5],loc[31][6],loc[31][7],loc[31][8],loc[31][9],loc[31][10]};end
            32:begin W21 = {loc[32][1],loc[32][2],loc[32][3],loc[32][4],loc[32][5],loc[32][6],loc[32][7],loc[32][8],loc[32][9],loc[32][10]};end
            33:begin W21 = {loc[33][1],loc[33][2],loc[33][3],loc[33][4],loc[33][5],loc[33][6],loc[33][7],loc[33][8],loc[33][9],loc[33][10]};end
            34:begin W21 = {loc[34][1],loc[34][2],loc[34][3],loc[34][4],loc[34][5],loc[34][6],loc[34][7],loc[34][8],loc[34][9],loc[34][10]};end
            35:begin W21 = {loc[35][1],loc[35][2],loc[35][3],loc[35][4],loc[35][5],loc[35][6],loc[35][7],loc[35][8],loc[35][9],loc[35][10]};end
            36:begin W21 = {loc[36][1],loc[36][2],loc[36][3],loc[36][4],loc[36][5],loc[36][6],loc[36][7],loc[36][8],loc[36][9],loc[36][10]};end
            37:begin W21 = {loc[37][1],loc[37][2],loc[37][3],loc[37][4],loc[37][5],loc[37][6],loc[37][7],loc[37][8],loc[37][9],loc[37][10]};end
            38:begin W21 = {loc[38][1],loc[38][2],loc[38][3],loc[38][4],loc[38][5],loc[38][6],loc[38][7],loc[38][8],loc[38][9],loc[38][10]};end
            39:begin W21 = {loc[39][1],loc[39][2],loc[39][3],loc[39][4],loc[39][5],loc[39][6],loc[39][7],loc[39][8],loc[39][9],loc[39][10]};end
            40:begin W21 = {loc[40][1],loc[40][2],loc[40][3],loc[40][4],loc[40][5],loc[40][6],loc[40][7],loc[40][8],loc[40][9],loc[40][10]};end
            41:begin W21 = {loc[41][1],loc[41][2],loc[41][3],loc[41][4],loc[41][5],loc[41][6],loc[41][7],loc[41][8],loc[41][9],loc[41][10]};end
            42:begin W21 = {loc[42][1],loc[42][2],loc[42][3],loc[42][4],loc[42][5],loc[42][6],loc[42][7],loc[42][8],loc[42][9],loc[42][10]};end
            43:begin W21 = {loc[43][1],loc[43][2],loc[43][3],loc[43][4],loc[43][5],loc[43][6],loc[43][7],loc[43][8],loc[43][9],loc[43][10]};end
            44:begin W21 = {loc[44][1],loc[44][2],loc[44][3],loc[44][4],loc[44][5],loc[44][6],loc[44][7],loc[44][8],loc[44][9],loc[44][10]};end
            45:begin W21 = {loc[45][1],loc[45][2],loc[45][3],loc[45][4],loc[45][5],loc[45][6],loc[45][7],loc[45][8],loc[45][9],loc[45][10]};end
            46:begin W21 = {loc[46][1],loc[46][2],loc[46][3],loc[46][4],loc[46][5],loc[46][6],loc[46][7],loc[46][8],loc[46][9],loc[46][10]};end
            47:begin W21 = {loc[47][1],loc[47][2],loc[47][3],loc[47][4],loc[47][5],loc[47][6],loc[47][7],loc[47][8],loc[47][9],loc[47][10]};end
            48:begin W21 = {loc[48][1],loc[48][2],loc[48][3],loc[48][4],loc[48][5],loc[48][6],loc[48][7],loc[48][8],loc[48][9],loc[48][10]};end
            49:begin W21 = {loc[49][1],loc[49][2],loc[49][3],loc[49][4],loc[49][5],loc[49][6],loc[49][7],loc[49][8],loc[49][9],loc[49][10]};end
            50:begin W21 = {loc[50][1],loc[50][2],loc[50][3],loc[50][4],loc[50][5],loc[50][6],loc[50][7],loc[50][8],loc[50][9],loc[50][10]};end
            51:begin W21 = {loc[51][1],loc[51][2],loc[51][3],loc[51][4],loc[51][5],loc[51][6],loc[51][7],loc[51][8],loc[51][9],loc[51][10]};end
            52:begin W21 = {loc[52][1],loc[52][2],loc[52][3],loc[52][4],loc[52][5],loc[52][6],loc[52][7],loc[52][8],loc[52][9],loc[52][10]};end
            53:begin W21 = {loc[53][1],loc[53][2],loc[53][3],loc[53][4],loc[53][5],loc[53][6],loc[53][7],loc[53][8],loc[53][9],loc[53][10]};end
            54:begin W21 = {loc[54][1],loc[54][2],loc[54][3],loc[54][4],loc[54][5],loc[54][6],loc[54][7],loc[54][8],loc[54][9],loc[54][10]};end
            55:begin W21 = {loc[55][1],loc[55][2],loc[55][3],loc[55][4],loc[55][5],loc[55][6],loc[55][7],loc[55][8],loc[55][9],loc[55][10]};end
            56:begin W21 = {loc[56][1],loc[56][2],loc[56][3],loc[56][4],loc[56][5],loc[56][6],loc[56][7],loc[56][8],loc[56][9],loc[56][10]};end
            57:begin W21 = {loc[57][1],loc[57][2],loc[57][3],loc[57][4],loc[57][5],loc[57][6],loc[57][7],loc[57][8],loc[57][9],loc[57][10]};end
            58:begin W21 = {loc[58][1],loc[58][2],loc[58][3],loc[58][4],loc[58][5],loc[58][6],loc[58][7],loc[58][8],loc[58][9],loc[58][10]};end
            59:begin W21 = {loc[59][1],loc[59][2],loc[59][3],loc[59][4],loc[59][5],loc[59][6],loc[59][7],loc[59][8],loc[59][9],loc[59][10]};end
            60:begin W21 = {loc[60][1],loc[60][2],loc[60][3],loc[60][4],loc[60][5],loc[60][6],loc[60][7],loc[60][8],loc[60][9],loc[60][10]};end
            61:begin W21 = {loc[61][1],loc[61][2],loc[61][3],loc[61][4],loc[61][5],loc[61][6],loc[61][7],loc[61][8],loc[61][9],loc[61][10]};end
            62:begin W21 = {loc[62][1],loc[62][2],loc[62][3],loc[62][4],loc[62][5],loc[62][6],loc[62][7],loc[62][8],loc[62][9],loc[62][10]};end
            63:begin W21 = {loc[63][1],loc[63][2],loc[63][3],loc[63][4],loc[63][5],loc[63][6],loc[63][7],loc[63][8],loc[63][9],loc[63][10]};end
            64:begin W21 = {loc[64][1],loc[64][2],loc[64][3],loc[64][4],loc[64][5],loc[64][6],loc[64][7],loc[64][8],loc[64][9],loc[64][10]};end
            65:begin W21 = {loc[65][1],loc[65][2],loc[65][3],loc[65][4],loc[65][5],loc[65][6],loc[65][7],loc[65][8],loc[65][9],loc[65][10]};end
            66:begin W21 = {loc[66][1],loc[66][2],loc[66][3],loc[66][4],loc[66][5],loc[66][6],loc[66][7],loc[66][8],loc[66][9],loc[66][10]};end
            67:begin W21 = {loc[67][1],loc[67][2],loc[67][3],loc[67][4],loc[67][5],loc[67][6],loc[67][7],loc[67][8],loc[67][9],loc[67][10]};end
            68:begin W21 = {loc[68][1],loc[68][2],loc[68][3],loc[68][4],loc[68][5],loc[68][6],loc[68][7],loc[68][8],loc[68][9],loc[68][10]};end
            69:begin W21 = {loc[69][1],loc[69][2],loc[69][3],loc[69][4],loc[69][5],loc[69][6],loc[69][7],loc[69][8],loc[69][9],loc[69][10]};end
            70:begin W21 = {loc[70][1],loc[70][2],loc[70][3],loc[70][4],loc[70][5],loc[70][6],loc[70][7],loc[70][8],loc[70][9],loc[70][10]};end
            71:begin W21 = {loc[71][1],loc[71][2],loc[71][3],loc[71][4],loc[71][5],loc[71][6],loc[71][7],loc[71][8],loc[71][9],loc[71][10]};end
            72:begin W21 = {loc[72][1],loc[72][2],loc[72][3],loc[72][4],loc[72][5],loc[72][6],loc[72][7],loc[72][8],loc[72][9],loc[72][10]};end
            73:begin W21 = {loc[73][1],loc[73][2],loc[73][3],loc[73][4],loc[73][5],loc[73][6],loc[73][7],loc[73][8],loc[73][9],loc[73][10]};end
            74:begin W21 = {loc[74][1],loc[74][2],loc[74][3],loc[74][4],loc[74][5],loc[74][6],loc[74][7],loc[74][8],loc[74][9],loc[74][10]};end
            75:begin W21 = {loc[75][1],loc[75][2],loc[75][3],loc[75][4],loc[75][5],loc[75][6],loc[75][7],loc[75][8],loc[75][9],loc[75][10]};end
            76:begin W21 = {loc[76][1],loc[76][2],loc[76][3],loc[76][4],loc[76][5],loc[76][6],loc[76][7],loc[76][8],loc[76][9],loc[76][10]};end
            77:begin W21 = {loc[77][1],loc[77][2],loc[77][3],loc[77][4],loc[77][5],loc[77][6],loc[77][7],loc[77][8],loc[77][9],loc[77][10]};end
            78:begin W21 = {loc[78][1],loc[78][2],loc[78][3],loc[78][4],loc[78][5],loc[78][6],loc[78][7],loc[78][8],loc[78][9],loc[78][10]};end
            79:begin W21 = {loc[79][1],loc[79][2],loc[79][3],loc[79][4],loc[79][5],loc[79][6],loc[79][7],loc[79][8],loc[79][9],loc[79][10]};end
            80:begin W21 = {loc[80][1],loc[80][2],loc[80][3],loc[80][4],loc[80][5],loc[80][6],loc[80][7],loc[80][8],loc[80][9],loc[80][10]};end
            81:begin W21 = {loc[81][1],loc[81][2],loc[81][3],loc[81][4],loc[81][5],loc[81][6],loc[81][7],loc[81][8],loc[81][9],loc[81][10]};end
            82:begin W21 = {loc[82][1],loc[82][2],loc[82][3],loc[82][4],loc[82][5],loc[82][6],loc[82][7],loc[82][8],loc[82][9],loc[82][10]};end
            83:begin W21 = {loc[83][1],loc[83][2],loc[83][3],loc[83][4],loc[83][5],loc[83][6],loc[83][7],loc[83][8],loc[83][9],loc[83][10]};end
            84:begin W21 = {loc[84][1],loc[84][2],loc[84][3],loc[84][4],loc[84][5],loc[84][6],loc[84][7],loc[84][8],loc[84][9],loc[84][10]};end
            85:begin W21 = {loc[85][1],loc[85][2],loc[85][3],loc[85][4],loc[85][5],loc[85][6],loc[85][7],loc[85][8],loc[85][9],loc[85][10]};end
            86:begin W21 = {loc[86][1],loc[86][2],loc[86][3],loc[86][4],loc[86][5],loc[86][6],loc[86][7],loc[86][8],loc[86][9],loc[86][10]};end
            87:begin W21 = {loc[87][1],loc[87][2],loc[87][3],loc[87][4],loc[87][5],loc[87][6],loc[87][7],loc[87][8],loc[87][9],loc[87][10]};end
            88:begin W21 = {loc[88][1],loc[88][2],loc[88][3],loc[88][4],loc[88][5],loc[88][6],loc[88][7],loc[88][8],loc[88][9],loc[88][10]};end
            89:begin W21 = {loc[89][1],loc[89][2],loc[89][3],loc[89][4],loc[89][5],loc[89][6],loc[89][7],loc[89][8],loc[89][9],loc[89][10]};end
            90:begin W21 = {loc[90][1],loc[90][2],loc[90][3],loc[90][4],loc[90][5],loc[90][6],loc[90][7],loc[90][8],loc[90][9],loc[90][10]};end
            91:begin W21 = {loc[91][1],loc[91][2],loc[91][3],loc[91][4],loc[91][5],loc[91][6],loc[91][7],loc[91][8],loc[91][9],loc[91][10]};end
            92:begin W21 = {loc[92][1],loc[92][2],loc[92][3],loc[92][4],loc[92][5],loc[92][6],loc[92][7],loc[92][8],loc[92][9],loc[92][10]};end
            93:begin W21 = {loc[93][1],loc[93][2],loc[93][3],loc[93][4],loc[93][5],loc[93][6],loc[93][7],loc[93][8],loc[93][9],loc[93][10]};end
            94:begin W21 = {loc[94][1],loc[94][2],loc[94][3],loc[94][4],loc[94][5],loc[94][6],loc[94][7],loc[94][8],loc[94][9],loc[94][10]};end
            95:begin W21 = {loc[95][1],loc[95][2],loc[95][3],loc[95][4],loc[95][5],loc[95][6],loc[95][7],loc[95][8],loc[95][9],loc[95][10]};end
            96:begin W21 = {loc[96][1],loc[96][2],loc[96][3],loc[96][4],loc[96][5],loc[96][6],loc[96][7],loc[96][8],loc[96][9],loc[96][10]};end
            97:begin W21 = {loc[97][1],loc[97][2],loc[97][3],loc[97][4],loc[97][5],loc[97][6],loc[97][7],loc[97][8],loc[97][9],loc[97][10]};end
            98:begin W21 = {loc[98][1],loc[98][2],loc[98][3],loc[98][4],loc[98][5],loc[98][6],loc[98][7],loc[98][8],loc[98][9],loc[98][10]};end
            99:begin W21 = {loc[99][1],loc[99][2],loc[99][3],loc[99][4],loc[99][5],loc[99][6],loc[99][7],loc[99][8],loc[99][9],loc[99][10]};end
            100:begin W21 = {loc[100][1],loc[100][2],loc[100][3],loc[100][4],loc[100][5],loc[100][6],loc[100][7],loc[100][8],loc[100][9],loc[100][10]};end
            101:begin W21 = {loc[101][1],loc[101][2],loc[101][3],loc[101][4],loc[101][5],loc[101][6],loc[101][7],loc[101][8],loc[101][9],loc[101][10]};end
            102:begin W21 = {loc[102][1],loc[102][2],loc[102][3],loc[102][4],loc[102][5],loc[102][6],loc[102][7],loc[102][8],loc[102][9],loc[102][10]};end
            103:begin W21 = {loc[103][1],loc[103][2],loc[103][3],loc[103][4],loc[103][5],loc[103][6],loc[103][7],loc[103][8],loc[103][9],loc[103][10]};end
            104:begin W21 = {loc[104][1],loc[104][2],loc[104][3],loc[104][4],loc[104][5],loc[104][6],loc[104][7],loc[104][8],loc[104][9],loc[104][10]};end
            105:begin W21 = {loc[105][1],loc[105][2],loc[105][3],loc[105][4],loc[105][5],loc[105][6],loc[105][7],loc[105][8],loc[105][9],loc[105][10]};end
            106:begin W21 = {loc[106][1],loc[106][2],loc[106][3],loc[106][4],loc[106][5],loc[106][6],loc[106][7],loc[106][8],loc[106][9],loc[106][10]};end
            107:begin W21 = {loc[107][1],loc[107][2],loc[107][3],loc[107][4],loc[107][5],loc[107][6],loc[107][7],loc[107][8],loc[107][9],loc[107][10]};end
            108:begin W21 = {loc[108][1],loc[108][2],loc[108][3],loc[108][4],loc[108][5],loc[108][6],loc[108][7],loc[108][8],loc[108][9],loc[108][10]};end
            109:begin W21 = {loc[109][1],loc[109][2],loc[109][3],loc[109][4],loc[109][5],loc[109][6],loc[109][7],loc[109][8],loc[109][9],loc[109][10]};end
            110:begin W21 = {loc[110][1],loc[110][2],loc[110][3],loc[110][4],loc[110][5],loc[110][6],loc[110][7],loc[110][8],loc[110][9],loc[110][10]};end
            111:begin W21 = {loc[111][1],loc[111][2],loc[111][3],loc[111][4],loc[111][5],loc[111][6],loc[111][7],loc[111][8],loc[111][9],loc[111][10]};end
            112:begin W21 = {loc[112][1],loc[112][2],loc[112][3],loc[112][4],loc[112][5],loc[112][6],loc[112][7],loc[112][8],loc[112][9],loc[112][10]};end
            113:begin W21 = {loc[113][1],loc[113][2],loc[113][3],loc[113][4],loc[113][5],loc[113][6],loc[113][7],loc[113][8],loc[113][9],loc[113][10]};end
            114:begin W21 = {loc[114][1],loc[114][2],loc[114][3],loc[114][4],loc[114][5],loc[114][6],loc[114][7],loc[114][8],loc[114][9],loc[114][10]};end
            115:begin W21 = {loc[115][1],loc[115][2],loc[115][3],loc[115][4],loc[115][5],loc[115][6],loc[115][7],loc[115][8],loc[115][9],loc[115][10]};end
            116:begin W21 = {loc[116][1],loc[116][2],loc[116][3],loc[116][4],loc[116][5],loc[116][6],loc[116][7],loc[116][8],loc[116][9],loc[116][10]};end
            117:begin W21 = {loc[117][1],loc[117][2],loc[117][3],loc[117][4],loc[117][5],loc[117][6],loc[117][7],loc[117][8],loc[117][9],loc[117][10]};end
            118:begin W21 = {loc[118][1],loc[118][2],loc[118][3],loc[118][4],loc[118][5],loc[118][6],loc[118][7],loc[118][8],loc[118][9],loc[118][10]};end
            119:begin W21 = {loc[119][1],loc[119][2],loc[119][3],loc[119][4],loc[119][5],loc[119][6],loc[119][7],loc[119][8],loc[119][9],loc[119][10]};end
            120:begin W21 = {loc[120][1],loc[120][2],loc[120][3],loc[120][4],loc[120][5],loc[120][6],loc[120][7],loc[120][8],loc[120][9],loc[120][10]};end
            121:begin W21 = {loc[121][1],loc[121][2],loc[121][3],loc[121][4],loc[121][5],loc[121][6],loc[121][7],loc[121][8],loc[121][9],loc[121][10]};end
            122:begin W21 = {loc[122][1],loc[122][2],loc[122][3],loc[122][4],loc[122][5],loc[122][6],loc[122][7],loc[122][8],loc[122][9],loc[122][10]};end
            123:begin W21 = {loc[123][1],loc[123][2],loc[123][3],loc[123][4],loc[123][5],loc[123][6],loc[123][7],loc[123][8],loc[123][9],loc[123][10]};end
            124:begin W21 = {loc[124][1],loc[124][2],loc[124][3],loc[124][4],loc[124][5],loc[124][6],loc[124][7],loc[124][8],loc[124][9],loc[124][10]};end
            125:begin W21 = {loc[125][1],loc[125][2],loc[125][3],loc[125][4],loc[125][5],loc[125][6],loc[125][7],loc[125][8],loc[125][9],loc[125][10]};end
            126:begin W21 = {loc[126][1],loc[126][2],loc[126][3],loc[126][4],loc[126][5],loc[126][6],loc[126][7],loc[126][8],loc[126][9],loc[126][10]};end
            127:begin W21 = {loc[127][1],loc[127][2],loc[127][3],loc[127][4],loc[127][5],loc[127][6],loc[127][7],loc[127][8],loc[127][9],loc[127][10]};end
            128:begin W21 = {loc[128][1],loc[128][2],loc[128][3],loc[128][4],loc[128][5],loc[128][6],loc[128][7],loc[128][8],loc[128][9],loc[128][10]};end
            129:begin W21 = {loc[129][1],loc[129][2],loc[129][3],loc[129][4],loc[129][5],loc[129][6],loc[129][7],loc[129][8],loc[129][9],loc[129][10]};end
            130:begin W21 = {loc[130][1],loc[130][2],loc[130][3],loc[130][4],loc[130][5],loc[130][6],loc[130][7],loc[130][8],loc[130][9],loc[130][10]};end
            131:begin W21 = {loc[131][1],loc[131][2],loc[131][3],loc[131][4],loc[131][5],loc[131][6],loc[131][7],loc[131][8],loc[131][9],loc[131][10]};end
            132:begin W21 = {loc[132][1],loc[132][2],loc[132][3],loc[132][4],loc[132][5],loc[132][6],loc[132][7],loc[132][8],loc[132][9],loc[132][10]};end
            133:begin W21 = {loc[133][1],loc[133][2],loc[133][3],loc[133][4],loc[133][5],loc[133][6],loc[133][7],loc[133][8],loc[133][9],loc[133][10]};end
            134:begin W21 = {loc[134][1],loc[134][2],loc[134][3],loc[134][4],loc[134][5],loc[134][6],loc[134][7],loc[134][8],loc[134][9],loc[134][10]};end
            135:begin W21 = {loc[135][1],loc[135][2],loc[135][3],loc[135][4],loc[135][5],loc[135][6],loc[135][7],loc[135][8],loc[135][9],loc[135][10]};end
            136:begin W21 = {loc[136][1],loc[136][2],loc[136][3],loc[136][4],loc[136][5],loc[136][6],loc[136][7],loc[136][8],loc[136][9],loc[136][10]};end
            137:begin W21 = {loc[137][1],loc[137][2],loc[137][3],loc[137][4],loc[137][5],loc[137][6],loc[137][7],loc[137][8],loc[137][9],loc[137][10]};end
            138:begin W21 = {loc[138][1],loc[138][2],loc[138][3],loc[138][4],loc[138][5],loc[138][6],loc[138][7],loc[138][8],loc[138][9],loc[138][10]};end
            139:begin W21 = {loc[139][1],loc[139][2],loc[139][3],loc[139][4],loc[139][5],loc[139][6],loc[139][7],loc[139][8],loc[139][9],loc[139][10]};end
            140:begin W21 = {loc[140][1],loc[140][2],loc[140][3],loc[140][4],loc[140][5],loc[140][6],loc[140][7],loc[140][8],loc[140][9],loc[140][10]};end
            141:begin W21 = {loc[141][1],loc[141][2],loc[141][3],loc[141][4],loc[141][5],loc[141][6],loc[141][7],loc[141][8],loc[141][9],loc[141][10]};end
            142:begin W21 = {loc[142][1],loc[142][2],loc[142][3],loc[142][4],loc[142][5],loc[142][6],loc[142][7],loc[142][8],loc[142][9],loc[142][10]};end
            143:begin W21 = {loc[143][1],loc[143][2],loc[143][3],loc[143][4],loc[143][5],loc[143][6],loc[143][7],loc[143][8],loc[143][9],loc[143][10]};end
            144:begin W21 = {loc[144][1],loc[144][2],loc[144][3],loc[144][4],loc[144][5],loc[144][6],loc[144][7],loc[144][8],loc[144][9],loc[144][10]};end
            145:begin W21 = {loc[145][1],loc[145][2],loc[145][3],loc[145][4],loc[145][5],loc[145][6],loc[145][7],loc[145][8],loc[145][9],loc[145][10]};end
            146:begin W21 = {loc[146][1],loc[146][2],loc[146][3],loc[146][4],loc[146][5],loc[146][6],loc[146][7],loc[146][8],loc[146][9],loc[146][10]};end
            147:begin W21 = {loc[147][1],loc[147][2],loc[147][3],loc[147][4],loc[147][5],loc[147][6],loc[147][7],loc[147][8],loc[147][9],loc[147][10]};end
            148:begin W21 = {loc[148][1],loc[148][2],loc[148][3],loc[148][4],loc[148][5],loc[148][6],loc[148][7],loc[148][8],loc[148][9],loc[148][10]};end
            149:begin W21 = {loc[149][1],loc[149][2],loc[149][3],loc[149][4],loc[149][5],loc[149][6],loc[149][7],loc[149][8],loc[149][9],loc[149][10]};end
            150:begin W21 = {loc[150][1],loc[150][2],loc[150][3],loc[150][4],loc[150][5],loc[150][6],loc[150][7],loc[150][8],loc[150][9],loc[150][10]};end
            151:begin W21 = {loc[151][1],loc[151][2],loc[151][3],loc[151][4],loc[151][5],loc[151][6],loc[151][7],loc[151][8],loc[151][9],loc[151][10]};end
            152:begin W21 = {loc[152][1],loc[152][2],loc[152][3],loc[152][4],loc[152][5],loc[152][6],loc[152][7],loc[152][8],loc[152][9],loc[152][10]};end
            153:begin W21 = {loc[153][1],loc[153][2],loc[153][3],loc[153][4],loc[153][5],loc[153][6],loc[153][7],loc[153][8],loc[153][9],loc[153][10]};end
            154:begin W21 = {loc[154][1],loc[154][2],loc[154][3],loc[154][4],loc[154][5],loc[154][6],loc[154][7],loc[154][8],loc[154][9],loc[154][10]};end
            155:begin W21 = {loc[155][1],loc[155][2],loc[155][3],loc[155][4],loc[155][5],loc[155][6],loc[155][7],loc[155][8],loc[155][9],loc[155][10]};end
            156:begin W21 = {loc[156][1],loc[156][2],loc[156][3],loc[156][4],loc[156][5],loc[156][6],loc[156][7],loc[156][8],loc[156][9],loc[156][10]};end
            157:begin W21 = {loc[157][1],loc[157][2],loc[157][3],loc[157][4],loc[157][5],loc[157][6],loc[157][7],loc[157][8],loc[157][9],loc[157][10]};end
            158:begin W21 = {loc[158][1],loc[158][2],loc[158][3],loc[158][4],loc[158][5],loc[158][6],loc[158][7],loc[158][8],loc[158][9],loc[158][10]};end
            159:begin W21 = {loc[159][1],loc[159][2],loc[159][3],loc[159][4],loc[159][5],loc[159][6],loc[159][7],loc[159][8],loc[159][9],loc[159][10]};end
            160:begin W21 = {loc[160][1],loc[160][2],loc[160][3],loc[160][4],loc[160][5],loc[160][6],loc[160][7],loc[160][8],loc[160][9],loc[160][10]};end
            161:begin W21 = {loc[161][1],loc[161][2],loc[161][3],loc[161][4],loc[161][5],loc[161][6],loc[161][7],loc[161][8],loc[161][9],loc[161][10]};end
            162:begin W21 = {loc[162][1],loc[162][2],loc[162][3],loc[162][4],loc[162][5],loc[162][6],loc[162][7],loc[162][8],loc[162][9],loc[162][10]};end
            163:begin W21 = {loc[163][1],loc[163][2],loc[163][3],loc[163][4],loc[163][5],loc[163][6],loc[163][7],loc[163][8],loc[163][9],loc[163][10]};end
            164:begin W21 = {loc[164][1],loc[164][2],loc[164][3],loc[164][4],loc[164][5],loc[164][6],loc[164][7],loc[164][8],loc[164][9],loc[164][10]};end
            165:begin W21 = {loc[165][1],loc[165][2],loc[165][3],loc[165][4],loc[165][5],loc[165][6],loc[165][7],loc[165][8],loc[165][9],loc[165][10]};end
            166:begin W21 = {loc[166][1],loc[166][2],loc[166][3],loc[166][4],loc[166][5],loc[166][6],loc[166][7],loc[166][8],loc[166][9],loc[166][10]};end
            167:begin W21 = {loc[167][1],loc[167][2],loc[167][3],loc[167][4],loc[167][5],loc[167][6],loc[167][7],loc[167][8],loc[167][9],loc[167][10]};end
            168:begin W21 = {loc[168][1],loc[168][2],loc[168][3],loc[168][4],loc[168][5],loc[168][6],loc[168][7],loc[168][8],loc[168][9],loc[168][10]};end
            169:begin W21 = {loc[169][1],loc[169][2],loc[169][3],loc[169][4],loc[169][5],loc[169][6],loc[169][7],loc[169][8],loc[169][9],loc[169][10]};end
            170:begin W21 = {loc[170][1],loc[170][2],loc[170][3],loc[170][4],loc[170][5],loc[170][6],loc[170][7],loc[170][8],loc[170][9],loc[170][10]};end
            171:begin W21 = {loc[171][1],loc[171][2],loc[171][3],loc[171][4],loc[171][5],loc[171][6],loc[171][7],loc[171][8],loc[171][9],loc[171][10]};end
            172:begin W21 = {loc[172][1],loc[172][2],loc[172][3],loc[172][4],loc[172][5],loc[172][6],loc[172][7],loc[172][8],loc[172][9],loc[172][10]};end
            173:begin W21 = {loc[173][1],loc[173][2],loc[173][3],loc[173][4],loc[173][5],loc[173][6],loc[173][7],loc[173][8],loc[173][9],loc[173][10]};end
            174:begin W21 = {loc[174][1],loc[174][2],loc[174][3],loc[174][4],loc[174][5],loc[174][6],loc[174][7],loc[174][8],loc[174][9],loc[174][10]};end
            175:begin W21 = {loc[175][1],loc[175][2],loc[175][3],loc[175][4],loc[175][5],loc[175][6],loc[175][7],loc[175][8],loc[175][9],loc[175][10]};end
            176:begin W21 = {loc[176][1],loc[176][2],loc[176][3],loc[176][4],loc[176][5],loc[176][6],loc[176][7],loc[176][8],loc[176][9],loc[176][10]};end
            177:begin W21 = {loc[177][1],loc[177][2],loc[177][3],loc[177][4],loc[177][5],loc[177][6],loc[177][7],loc[177][8],loc[177][9],loc[177][10]};end
            178:begin W21 = {loc[178][1],loc[178][2],loc[178][3],loc[178][4],loc[178][5],loc[178][6],loc[178][7],loc[178][8],loc[178][9],loc[178][10]};end
            179:begin W21 = {loc[179][1],loc[179][2],loc[179][3],loc[179][4],loc[179][5],loc[179][6],loc[179][7],loc[179][8],loc[179][9],loc[179][10]};end
            180:begin W21 = {loc[180][1],loc[180][2],loc[180][3],loc[180][4],loc[180][5],loc[180][6],loc[180][7],loc[180][8],loc[180][9],loc[180][10]};end
            181:begin W21 = {loc[181][1],loc[181][2],loc[181][3],loc[181][4],loc[181][5],loc[181][6],loc[181][7],loc[181][8],loc[181][9],loc[181][10]};end
            182:begin W21 = {loc[182][1],loc[182][2],loc[182][3],loc[182][4],loc[182][5],loc[182][6],loc[182][7],loc[182][8],loc[182][9],loc[182][10]};end
            183:begin W21 = {loc[183][1],loc[183][2],loc[183][3],loc[183][4],loc[183][5],loc[183][6],loc[183][7],loc[183][8],loc[183][9],loc[183][10]};end
            184:begin W21 = {loc[184][1],loc[184][2],loc[184][3],loc[184][4],loc[184][5],loc[184][6],loc[184][7],loc[184][8],loc[184][9],loc[184][10]};end
            185:begin W21 = {loc[185][1],loc[185][2],loc[185][3],loc[185][4],loc[185][5],loc[185][6],loc[185][7],loc[185][8],loc[185][9],loc[185][10]};end
            186:begin W21 = {loc[186][1],loc[186][2],loc[186][3],loc[186][4],loc[186][5],loc[186][6],loc[186][7],loc[186][8],loc[186][9],loc[186][10]};end
            187:begin W21 = {loc[187][1],loc[187][2],loc[187][3],loc[187][4],loc[187][5],loc[187][6],loc[187][7],loc[187][8],loc[187][9],loc[187][10]};end
            188:begin W21 = {loc[188][1],loc[188][2],loc[188][3],loc[188][4],loc[188][5],loc[188][6],loc[188][7],loc[188][8],loc[188][9],loc[188][10]};end
            189:begin W21 = {loc[189][1],loc[189][2],loc[189][3],loc[189][4],loc[189][5],loc[189][6],loc[189][7],loc[189][8],loc[189][9],loc[189][10]};end
            190:begin W21 = {loc[190][1],loc[190][2],loc[190][3],loc[190][4],loc[190][5],loc[190][6],loc[190][7],loc[190][8],loc[190][9],loc[190][10]};end
            191:begin W21 = {loc[191][1],loc[191][2],loc[191][3],loc[191][4],loc[191][5],loc[191][6],loc[191][7],loc[191][8],loc[191][9],loc[191][10]};end
            192:begin W21 = {loc[192][1],loc[192][2],loc[192][3],loc[192][4],loc[192][5],loc[192][6],loc[192][7],loc[192][8],loc[192][9],loc[192][10]};end
            193:begin W21 = {loc[193][1],loc[193][2],loc[193][3],loc[193][4],loc[193][5],loc[193][6],loc[193][7],loc[193][8],loc[193][9],loc[193][10]};end
            194:begin W21 = {loc[194][1],loc[194][2],loc[194][3],loc[194][4],loc[194][5],loc[194][6],loc[194][7],loc[194][8],loc[194][9],loc[194][10]};end
            195:begin W21 = {loc[195][1],loc[195][2],loc[195][3],loc[195][4],loc[195][5],loc[195][6],loc[195][7],loc[195][8],loc[195][9],loc[195][10]};end
            196:begin W21 = {loc[196][1],loc[196][2],loc[196][3],loc[196][4],loc[196][5],loc[196][6],loc[196][7],loc[196][8],loc[196][9],loc[196][10]};end
            197:begin W21 = {loc[197][1],loc[197][2],loc[197][3],loc[197][4],loc[197][5],loc[197][6],loc[197][7],loc[197][8],loc[197][9],loc[197][10]};end
            198:begin W21 = {loc[198][1],loc[198][2],loc[198][3],loc[198][4],loc[198][5],loc[198][6],loc[198][7],loc[198][8],loc[198][9],loc[198][10]};end
            199:begin W21 = {loc[199][1],loc[199][2],loc[199][3],loc[199][4],loc[199][5],loc[199][6],loc[199][7],loc[199][8],loc[199][9],loc[199][10]};end
            200:begin W21 = {loc[200][1],loc[200][2],loc[200][3],loc[200][4],loc[200][5],loc[200][6],loc[200][7],loc[200][8],loc[200][9],loc[200][10]};end
            201:begin W21 = {loc[201][1],loc[201][2],loc[201][3],loc[201][4],loc[201][5],loc[201][6],loc[201][7],loc[201][8],loc[201][9],loc[201][10]};end
            202:begin W21 = {loc[202][1],loc[202][2],loc[202][3],loc[202][4],loc[202][5],loc[202][6],loc[202][7],loc[202][8],loc[202][9],loc[202][10]};end
            203:begin W21 = {loc[203][1],loc[203][2],loc[203][3],loc[203][4],loc[203][5],loc[203][6],loc[203][7],loc[203][8],loc[203][9],loc[203][10]};end
            204:begin W21 = {loc[204][1],loc[204][2],loc[204][3],loc[204][4],loc[204][5],loc[204][6],loc[204][7],loc[204][8],loc[204][9],loc[204][10]};end
            205:begin W21 = {loc[205][1],loc[205][2],loc[205][3],loc[205][4],loc[205][5],loc[205][6],loc[205][7],loc[205][8],loc[205][9],loc[205][10]};end
            206:begin W21 = {loc[206][1],loc[206][2],loc[206][3],loc[206][4],loc[206][5],loc[206][6],loc[206][7],loc[206][8],loc[206][9],loc[206][10]};end
            207:begin W21 = {loc[207][1],loc[207][2],loc[207][3],loc[207][4],loc[207][5],loc[207][6],loc[207][7],loc[207][8],loc[207][9],loc[207][10]};end
            208:begin W21 = {loc[208][1],loc[208][2],loc[208][3],loc[208][4],loc[208][5],loc[208][6],loc[208][7],loc[208][8],loc[208][9],loc[208][10]};end
            209:begin W21 = {loc[209][1],loc[209][2],loc[209][3],loc[209][4],loc[209][5],loc[209][6],loc[209][7],loc[209][8],loc[209][9],loc[209][10]};end
            210:begin W21 = {loc[210][1],loc[210][2],loc[210][3],loc[210][4],loc[210][5],loc[210][6],loc[210][7],loc[210][8],loc[210][9],loc[210][10]};end
            211:begin W21 = {loc[211][1],loc[211][2],loc[211][3],loc[211][4],loc[211][5],loc[211][6],loc[211][7],loc[211][8],loc[211][9],loc[211][10]};end
            212:begin W21 = {loc[212][1],loc[212][2],loc[212][3],loc[212][4],loc[212][5],loc[212][6],loc[212][7],loc[212][8],loc[212][9],loc[212][10]};end
            213:begin W21 = {loc[213][1],loc[213][2],loc[213][3],loc[213][4],loc[213][5],loc[213][6],loc[213][7],loc[213][8],loc[213][9],loc[213][10]};end
            214:begin W21 = {loc[214][1],loc[214][2],loc[214][3],loc[214][4],loc[214][5],loc[214][6],loc[214][7],loc[214][8],loc[214][9],loc[214][10]};end
            215:begin W21 = {loc[215][1],loc[215][2],loc[215][3],loc[215][4],loc[215][5],loc[215][6],loc[215][7],loc[215][8],loc[215][9],loc[215][10]};end
            216:begin W21 = {loc[216][1],loc[216][2],loc[216][3],loc[216][4],loc[216][5],loc[216][6],loc[216][7],loc[216][8],loc[216][9],loc[216][10]};end
            217:begin W21 = {loc[217][1],loc[217][2],loc[217][3],loc[217][4],loc[217][5],loc[217][6],loc[217][7],loc[217][8],loc[217][9],loc[217][10]};end
            218:begin W21 = {loc[218][1],loc[218][2],loc[218][3],loc[218][4],loc[218][5],loc[218][6],loc[218][7],loc[218][8],loc[218][9],loc[218][10]};end
            219:begin W21 = {loc[219][1],loc[219][2],loc[219][3],loc[219][4],loc[219][5],loc[219][6],loc[219][7],loc[219][8],loc[219][9],loc[219][10]};end
            220:begin W21 = {loc[220][1],loc[220][2],loc[220][3],loc[220][4],loc[220][5],loc[220][6],loc[220][7],loc[220][8],loc[220][9],loc[220][10]};end
            221:begin W21 = {loc[221][1],loc[221][2],loc[221][3],loc[221][4],loc[221][5],loc[221][6],loc[221][7],loc[221][8],loc[221][9],loc[221][10]};end
            222:begin W21 = {loc[222][1],loc[222][2],loc[222][3],loc[222][4],loc[222][5],loc[222][6],loc[222][7],loc[222][8],loc[222][9],loc[222][10]};end
            223:begin W21 = {loc[223][1],loc[223][2],loc[223][3],loc[223][4],loc[223][5],loc[223][6],loc[223][7],loc[223][8],loc[223][9],loc[223][10]};end
            224:begin W21 = {loc[224][1],loc[224][2],loc[224][3],loc[224][4],loc[224][5],loc[224][6],loc[224][7],loc[224][8],loc[224][9],loc[224][10]};end
            225:begin W21 = {loc[225][1],loc[225][2],loc[225][3],loc[225][4],loc[225][5],loc[225][6],loc[225][7],loc[225][8],loc[225][9],loc[225][10]};end
            226:begin W21 = {loc[226][1],loc[226][2],loc[226][3],loc[226][4],loc[226][5],loc[226][6],loc[226][7],loc[226][8],loc[226][9],loc[226][10]};end
            227:begin W21 = {loc[227][1],loc[227][2],loc[227][3],loc[227][4],loc[227][5],loc[227][6],loc[227][7],loc[227][8],loc[227][9],loc[227][10]};end
            228:begin W21 = {loc[228][1],loc[228][2],loc[228][3],loc[228][4],loc[228][5],loc[228][6],loc[228][7],loc[228][8],loc[228][9],loc[228][10]};end
            229:begin W21 = {loc[229][1],loc[229][2],loc[229][3],loc[229][4],loc[229][5],loc[229][6],loc[229][7],loc[229][8],loc[229][9],loc[229][10]};end
            230:begin W21 = {loc[230][1],loc[230][2],loc[230][3],loc[230][4],loc[230][5],loc[230][6],loc[230][7],loc[230][8],loc[230][9],loc[230][10]};end
            231:begin W21 = {loc[231][1],loc[231][2],loc[231][3],loc[231][4],loc[231][5],loc[231][6],loc[231][7],loc[231][8],loc[231][9],loc[231][10]};end
            232:begin W21 = {loc[232][1],loc[232][2],loc[232][3],loc[232][4],loc[232][5],loc[232][6],loc[232][7],loc[232][8],loc[232][9],loc[232][10]};end
            233:begin W21 = {loc[233][1],loc[233][2],loc[233][3],loc[233][4],loc[233][5],loc[233][6],loc[233][7],loc[233][8],loc[233][9],loc[233][10]};end
            234:begin W21 = {loc[234][1],loc[234][2],loc[234][3],loc[234][4],loc[234][5],loc[234][6],loc[234][7],loc[234][8],loc[234][9],loc[234][10]};end
            235:begin W21 = {loc[235][1],loc[235][2],loc[235][3],loc[235][4],loc[235][5],loc[235][6],loc[235][7],loc[235][8],loc[235][9],loc[235][10]};end
            236:begin W21 = {loc[236][1],loc[236][2],loc[236][3],loc[236][4],loc[236][5],loc[236][6],loc[236][7],loc[236][8],loc[236][9],loc[236][10]};end
            237:begin W21 = {loc[237][1],loc[237][2],loc[237][3],loc[237][4],loc[237][5],loc[237][6],loc[237][7],loc[237][8],loc[237][9],loc[237][10]};end
            238:begin W21 = {loc[238][1],loc[238][2],loc[238][3],loc[238][4],loc[238][5],loc[238][6],loc[238][7],loc[238][8],loc[238][9],loc[238][10]};end
            239:begin W21 = {loc[239][1],loc[239][2],loc[239][3],loc[239][4],loc[239][5],loc[239][6],loc[239][7],loc[239][8],loc[239][9],loc[239][10]};end
            240:begin W21 = {loc[240][1],loc[240][2],loc[240][3],loc[240][4],loc[240][5],loc[240][6],loc[240][7],loc[240][8],loc[240][9],loc[240][10]};end
            241:begin W21 = {loc[241][1],loc[241][2],loc[241][3],loc[241][4],loc[241][5],loc[241][6],loc[241][7],loc[241][8],loc[241][9],loc[241][10]};end
            242:begin W21 = {loc[242][1],loc[242][2],loc[242][3],loc[242][4],loc[242][5],loc[242][6],loc[242][7],loc[242][8],loc[242][9],loc[242][10]};end
            243:begin W21 = {loc[243][1],loc[243][2],loc[243][3],loc[243][4],loc[243][5],loc[243][6],loc[243][7],loc[243][8],loc[243][9],loc[243][10]};end
            244:begin W21 = {loc[244][1],loc[244][2],loc[244][3],loc[244][4],loc[244][5],loc[244][6],loc[244][7],loc[244][8],loc[244][9],loc[244][10]};end
            245:begin W21 = {loc[245][1],loc[245][2],loc[245][3],loc[245][4],loc[245][5],loc[245][6],loc[245][7],loc[245][8],loc[245][9],loc[245][10]};end
            246:begin W21 = {loc[246][1],loc[246][2],loc[246][3],loc[246][4],loc[246][5],loc[246][6],loc[246][7],loc[246][8],loc[246][9],loc[246][10]};end
            247:begin W21 = {loc[247][1],loc[247][2],loc[247][3],loc[247][4],loc[247][5],loc[247][6],loc[247][7],loc[247][8],loc[247][9],loc[247][10]};end
            248:begin W21 = {loc[248][1],loc[248][2],loc[248][3],loc[248][4],loc[248][5],loc[248][6],loc[248][7],loc[248][8],loc[248][9],loc[248][10]};end
            249:begin W21 = {loc[249][1],loc[249][2],loc[249][3],loc[249][4],loc[249][5],loc[249][6],loc[249][7],loc[249][8],loc[249][9],loc[249][10]};end
            250:begin W21 = {loc[250][1],loc[250][2],loc[250][3],loc[250][4],loc[250][5],loc[250][6],loc[250][7],loc[250][8],loc[250][9],loc[250][10]};end
            251:begin W21 = {loc[251][1],loc[251][2],loc[251][3],loc[251][4],loc[251][5],loc[251][6],loc[251][7],loc[251][8],loc[251][9],loc[251][10]};end
            252:begin W21 = {loc[252][1],loc[252][2],loc[252][3],loc[252][4],loc[252][5],loc[252][6],loc[252][7],loc[252][8],loc[252][9],loc[252][10]};end
            253:begin W21 = {loc[253][1],loc[253][2],loc[253][3],loc[253][4],loc[253][5],loc[253][6],loc[253][7],loc[253][8],loc[253][9],loc[253][10]};end
            254:begin W21 = {loc[254][1],loc[254][2],loc[254][3],loc[254][4],loc[254][5],loc[254][6],loc[254][7],loc[254][8],loc[254][9],loc[254][10]};end
            255:begin W21 = {loc[255][1],loc[255][2],loc[255][3],loc[255][4],loc[255][5],loc[255][6],loc[255][7],loc[255][8],loc[255][9],loc[255][10]};end
            256:begin W21 = {loc[256][1],loc[256][2],loc[256][3],loc[256][4],loc[256][5],loc[256][6],loc[256][7],loc[256][8],loc[256][9],loc[256][10]};end
            257:begin W21 = {loc[257][1],loc[257][2],loc[257][3],loc[257][4],loc[257][5],loc[257][6],loc[257][7],loc[257][8],loc[257][9],loc[257][10]};end
            258:begin W21 = {loc[258][1],loc[258][2],loc[258][3],loc[258][4],loc[258][5],loc[258][6],loc[258][7],loc[258][8],loc[258][9],loc[258][10]};end
            259:begin W21 = {loc[259][1],loc[259][2],loc[259][3],loc[259][4],loc[259][5],loc[259][6],loc[259][7],loc[259][8],loc[259][9],loc[259][10]};end
            260:begin W21 = {loc[260][1],loc[260][2],loc[260][3],loc[260][4],loc[260][5],loc[260][6],loc[260][7],loc[260][8],loc[260][9],loc[260][10]};end
            261:begin W21 = {loc[261][1],loc[261][2],loc[261][3],loc[261][4],loc[261][5],loc[261][6],loc[261][7],loc[261][8],loc[261][9],loc[261][10]};end
            262:begin W21 = {loc[262][1],loc[262][2],loc[262][3],loc[262][4],loc[262][5],loc[262][6],loc[262][7],loc[262][8],loc[262][9],loc[262][10]};end
            263:begin W21 = {loc[263][1],loc[263][2],loc[263][3],loc[263][4],loc[263][5],loc[263][6],loc[263][7],loc[263][8],loc[263][9],loc[263][10]};end
            264:begin W21 = {loc[264][1],loc[264][2],loc[264][3],loc[264][4],loc[264][5],loc[264][6],loc[264][7],loc[264][8],loc[264][9],loc[264][10]};end
            265:begin W21 = {loc[265][1],loc[265][2],loc[265][3],loc[265][4],loc[265][5],loc[265][6],loc[265][7],loc[265][8],loc[265][9],loc[265][10]};end
            266:begin W21 = {loc[266][1],loc[266][2],loc[266][3],loc[266][4],loc[266][5],loc[266][6],loc[266][7],loc[266][8],loc[266][9],loc[266][10]};end
            267:begin W21 = {loc[267][1],loc[267][2],loc[267][3],loc[267][4],loc[267][5],loc[267][6],loc[267][7],loc[267][8],loc[267][9],loc[267][10]};end
            268:begin W21 = {loc[268][1],loc[268][2],loc[268][3],loc[268][4],loc[268][5],loc[268][6],loc[268][7],loc[268][8],loc[268][9],loc[268][10]};end
            269:begin W21 = {loc[269][1],loc[269][2],loc[269][3],loc[269][4],loc[269][5],loc[269][6],loc[269][7],loc[269][8],loc[269][9],loc[269][10]};end
            270:begin W21 = {loc[270][1],loc[270][2],loc[270][3],loc[270][4],loc[270][5],loc[270][6],loc[270][7],loc[270][8],loc[270][9],loc[270][10]};end
            271:begin W21 = {loc[271][1],loc[271][2],loc[271][3],loc[271][4],loc[271][5],loc[271][6],loc[271][7],loc[271][8],loc[271][9],loc[271][10]};end
            272:begin W21 = {loc[272][1],loc[272][2],loc[272][3],loc[272][4],loc[272][5],loc[272][6],loc[272][7],loc[272][8],loc[272][9],loc[272][10]};end
            273:begin W21 = {loc[273][1],loc[273][2],loc[273][3],loc[273][4],loc[273][5],loc[273][6],loc[273][7],loc[273][8],loc[273][9],loc[273][10]};end
            274:begin W21 = {loc[274][1],loc[274][2],loc[274][3],loc[274][4],loc[274][5],loc[274][6],loc[274][7],loc[274][8],loc[274][9],loc[274][10]};end
            275:begin W21 = {loc[275][1],loc[275][2],loc[275][3],loc[275][4],loc[275][5],loc[275][6],loc[275][7],loc[275][8],loc[275][9],loc[275][10]};end
            276:begin W21 = {loc[276][1],loc[276][2],loc[276][3],loc[276][4],loc[276][5],loc[276][6],loc[276][7],loc[276][8],loc[276][9],loc[276][10]};end
            277:begin W21 = {loc[277][1],loc[277][2],loc[277][3],loc[277][4],loc[277][5],loc[277][6],loc[277][7],loc[277][8],loc[277][9],loc[277][10]};end
            278:begin W21 = {loc[278][1],loc[278][2],loc[278][3],loc[278][4],loc[278][5],loc[278][6],loc[278][7],loc[278][8],loc[278][9],loc[278][10]};end
            279:begin W21 = {loc[279][1],loc[279][2],loc[279][3],loc[279][4],loc[279][5],loc[279][6],loc[279][7],loc[279][8],loc[279][9],loc[279][10]};end
            280:begin W21 = {loc[280][1],loc[280][2],loc[280][3],loc[280][4],loc[280][5],loc[280][6],loc[280][7],loc[280][8],loc[280][9],loc[280][10]};end
            281:begin W21 = {loc[281][1],loc[281][2],loc[281][3],loc[281][4],loc[281][5],loc[281][6],loc[281][7],loc[281][8],loc[281][9],loc[281][10]};end
            282:begin W21 = {loc[282][1],loc[282][2],loc[282][3],loc[282][4],loc[282][5],loc[282][6],loc[282][7],loc[282][8],loc[282][9],loc[282][10]};end
            283:begin W21 = {loc[283][1],loc[283][2],loc[283][3],loc[283][4],loc[283][5],loc[283][6],loc[283][7],loc[283][8],loc[283][9],loc[283][10]};end
            284:begin W21 = {loc[284][1],loc[284][2],loc[284][3],loc[284][4],loc[284][5],loc[284][6],loc[284][7],loc[284][8],loc[284][9],loc[284][10]};end
            285:begin W21 = {loc[285][1],loc[285][2],loc[285][3],loc[285][4],loc[285][5],loc[285][6],loc[285][7],loc[285][8],loc[285][9],loc[285][10]};end
            286:begin W21 = {loc[286][1],loc[286][2],loc[286][3],loc[286][4],loc[286][5],loc[286][6],loc[286][7],loc[286][8],loc[286][9],loc[286][10]};end
            287:begin W21 = {loc[287][1],loc[287][2],loc[287][3],loc[287][4],loc[287][5],loc[287][6],loc[287][7],loc[287][8],loc[287][9],loc[287][10]};end
            288:begin W21 = {loc[288][1],loc[288][2],loc[288][3],loc[288][4],loc[288][5],loc[288][6],loc[288][7],loc[288][8],loc[288][9],loc[288][10]};end
            289:begin W21 = {loc[289][1],loc[289][2],loc[289][3],loc[289][4],loc[289][5],loc[289][6],loc[289][7],loc[289][8],loc[289][9],loc[289][10]};end
            290:begin W21 = {loc[290][1],loc[290][2],loc[290][3],loc[290][4],loc[290][5],loc[290][6],loc[290][7],loc[290][8],loc[290][9],loc[290][10]};end
            291:begin W21 = {loc[291][1],loc[291][2],loc[291][3],loc[291][4],loc[291][5],loc[291][6],loc[291][7],loc[291][8],loc[291][9],loc[291][10]};end
            292:begin W21 = {loc[292][1],loc[292][2],loc[292][3],loc[292][4],loc[292][5],loc[292][6],loc[292][7],loc[292][8],loc[292][9],loc[292][10]};end
            293:begin W21 = {loc[293][1],loc[293][2],loc[293][3],loc[293][4],loc[293][5],loc[293][6],loc[293][7],loc[293][8],loc[293][9],loc[293][10]};end
            294:begin W21 = {loc[294][1],loc[294][2],loc[294][3],loc[294][4],loc[294][5],loc[294][6],loc[294][7],loc[294][8],loc[294][9],loc[294][10]};end
            295:begin W21 = {loc[295][1],loc[295][2],loc[295][3],loc[295][4],loc[295][5],loc[295][6],loc[295][7],loc[295][8],loc[295][9],loc[295][10]};end
            296:begin W21 = {loc[296][1],loc[296][2],loc[296][3],loc[296][4],loc[296][5],loc[296][6],loc[296][7],loc[296][8],loc[296][9],loc[296][10]};end
            297:begin W21 = {loc[297][1],loc[297][2],loc[297][3],loc[297][4],loc[297][5],loc[297][6],loc[297][7],loc[297][8],loc[297][9],loc[297][10]};end
            298:begin W21 = {loc[298][1],loc[298][2],loc[298][3],loc[298][4],loc[298][5],loc[298][6],loc[298][7],loc[298][8],loc[298][9],loc[298][10]};end
            299:begin W21 = {loc[299][1],loc[299][2],loc[299][3],loc[299][4],loc[299][5],loc[299][6],loc[299][7],loc[299][8],loc[299][9],loc[299][10]};end
            300:begin W21 = {loc[300][1],loc[300][2],loc[300][3],loc[300][4],loc[300][5],loc[300][6],loc[300][7],loc[300][8],loc[300][9],loc[300][10]};end
            301:begin W21 = {loc[301][1],loc[301][2],loc[301][3],loc[301][4],loc[301][5],loc[301][6],loc[301][7],loc[301][8],loc[301][9],loc[301][10]};end
            302:begin W21 = {loc[302][1],loc[302][2],loc[302][3],loc[302][4],loc[302][5],loc[302][6],loc[302][7],loc[302][8],loc[302][9],loc[302][10]};end
            303:begin W21 = {loc[303][1],loc[303][2],loc[303][3],loc[303][4],loc[303][5],loc[303][6],loc[303][7],loc[303][8],loc[303][9],loc[303][10]};end
            304:begin W21 = {loc[304][1],loc[304][2],loc[304][3],loc[304][4],loc[304][5],loc[304][6],loc[304][7],loc[304][8],loc[304][9],loc[304][10]};end
            305:begin W21 = {loc[305][1],loc[305][2],loc[305][3],loc[305][4],loc[305][5],loc[305][6],loc[305][7],loc[305][8],loc[305][9],loc[305][10]};end
            306:begin W21 = {loc[306][1],loc[306][2],loc[306][3],loc[306][4],loc[306][5],loc[306][6],loc[306][7],loc[306][8],loc[306][9],loc[306][10]};end
            307:begin W21 = {loc[307][1],loc[307][2],loc[307][3],loc[307][4],loc[307][5],loc[307][6],loc[307][7],loc[307][8],loc[307][9],loc[307][10]};end
            308:begin W21 = {loc[308][1],loc[308][2],loc[308][3],loc[308][4],loc[308][5],loc[308][6],loc[308][7],loc[308][8],loc[308][9],loc[308][10]};end
            309:begin W21 = {loc[309][1],loc[309][2],loc[309][3],loc[309][4],loc[309][5],loc[309][6],loc[309][7],loc[309][8],loc[309][9],loc[309][10]};end
            310:begin W21 = {loc[310][1],loc[310][2],loc[310][3],loc[310][4],loc[310][5],loc[310][6],loc[310][7],loc[310][8],loc[310][9],loc[310][10]};end
            311:begin W21 = {loc[311][1],loc[311][2],loc[311][3],loc[311][4],loc[311][5],loc[311][6],loc[311][7],loc[311][8],loc[311][9],loc[311][10]};end
            312:begin W21 = {loc[312][1],loc[312][2],loc[312][3],loc[312][4],loc[312][5],loc[312][6],loc[312][7],loc[312][8],loc[312][9],loc[312][10]};end
            313:begin W21 = {loc[313][1],loc[313][2],loc[313][3],loc[313][4],loc[313][5],loc[313][6],loc[313][7],loc[313][8],loc[313][9],loc[313][10]};end
            314:begin W21 = {loc[314][1],loc[314][2],loc[314][3],loc[314][4],loc[314][5],loc[314][6],loc[314][7],loc[314][8],loc[314][9],loc[314][10]};end
            315:begin W21 = {loc[315][1],loc[315][2],loc[315][3],loc[315][4],loc[315][5],loc[315][6],loc[315][7],loc[315][8],loc[315][9],loc[315][10]};end
            316:begin W21 = {loc[316][1],loc[316][2],loc[316][3],loc[316][4],loc[316][5],loc[316][6],loc[316][7],loc[316][8],loc[316][9],loc[316][10]};end
            317:begin W21 = {loc[317][1],loc[317][2],loc[317][3],loc[317][4],loc[317][5],loc[317][6],loc[317][7],loc[317][8],loc[317][9],loc[317][10]};end
            318:begin W21 = {loc[318][1],loc[318][2],loc[318][3],loc[318][4],loc[318][5],loc[318][6],loc[318][7],loc[318][8],loc[318][9],loc[318][10]};end
            319:begin W21 = {loc[319][1],loc[319][2],loc[319][3],loc[319][4],loc[319][5],loc[319][6],loc[319][7],loc[319][8],loc[319][9],loc[319][10]};end
            320:begin W21 = {loc[320][1],loc[320][2],loc[320][3],loc[320][4],loc[320][5],loc[320][6],loc[320][7],loc[320][8],loc[320][9],loc[320][10]};end
            321:begin W21 = {loc[321][1],loc[321][2],loc[321][3],loc[321][4],loc[321][5],loc[321][6],loc[321][7],loc[321][8],loc[321][9],loc[321][10]};end
            322:begin W21 = {loc[322][1],loc[322][2],loc[322][3],loc[322][4],loc[322][5],loc[322][6],loc[322][7],loc[322][8],loc[322][9],loc[322][10]};end
            323:begin W21 = {loc[323][1],loc[323][2],loc[323][3],loc[323][4],loc[323][5],loc[323][6],loc[323][7],loc[323][8],loc[323][9],loc[323][10]};end
            324:begin W21 = {loc[324][1],loc[324][2],loc[324][3],loc[324][4],loc[324][5],loc[324][6],loc[324][7],loc[324][8],loc[324][9],loc[324][10]};end
            325:begin W21 = {loc[325][1],loc[325][2],loc[325][3],loc[325][4],loc[325][5],loc[325][6],loc[325][7],loc[325][8],loc[325][9],loc[325][10]};end
            326:begin W21 = {loc[326][1],loc[326][2],loc[326][3],loc[326][4],loc[326][5],loc[326][6],loc[326][7],loc[326][8],loc[326][9],loc[326][10]};end
            327:begin W21 = {loc[327][1],loc[327][2],loc[327][3],loc[327][4],loc[327][5],loc[327][6],loc[327][7],loc[327][8],loc[327][9],loc[327][10]};end
            328:begin W21 = {loc[328][1],loc[328][2],loc[328][3],loc[328][4],loc[328][5],loc[328][6],loc[328][7],loc[328][8],loc[328][9],loc[328][10]};end
            329:begin W21 = {loc[329][1],loc[329][2],loc[329][3],loc[329][4],loc[329][5],loc[329][6],loc[329][7],loc[329][8],loc[329][9],loc[329][10]};end
            330:begin W21 = {loc[330][1],loc[330][2],loc[330][3],loc[330][4],loc[330][5],loc[330][6],loc[330][7],loc[330][8],loc[330][9],loc[330][10]};end
            331:begin W21 = {loc[331][1],loc[331][2],loc[331][3],loc[331][4],loc[331][5],loc[331][6],loc[331][7],loc[331][8],loc[331][9],loc[331][10]};end
            332:begin W21 = {loc[332][1],loc[332][2],loc[332][3],loc[332][4],loc[332][5],loc[332][6],loc[332][7],loc[332][8],loc[332][9],loc[332][10]};end
            333:begin W21 = {loc[333][1],loc[333][2],loc[333][3],loc[333][4],loc[333][5],loc[333][6],loc[333][7],loc[333][8],loc[333][9],loc[333][10]};end
            334:begin W21 = {loc[334][1],loc[334][2],loc[334][3],loc[334][4],loc[334][5],loc[334][6],loc[334][7],loc[334][8],loc[334][9],loc[334][10]};end
            335:begin W21 = {loc[335][1],loc[335][2],loc[335][3],loc[335][4],loc[335][5],loc[335][6],loc[335][7],loc[335][8],loc[335][9],loc[335][10]};end
            336:begin W21 = {loc[336][1],loc[336][2],loc[336][3],loc[336][4],loc[336][5],loc[336][6],loc[336][7],loc[336][8],loc[336][9],loc[336][10]};end
            337:begin W21 = {loc[337][1],loc[337][2],loc[337][3],loc[337][4],loc[337][5],loc[337][6],loc[337][7],loc[337][8],loc[337][9],loc[337][10]};end
            338:begin W21 = {loc[338][1],loc[338][2],loc[338][3],loc[338][4],loc[338][5],loc[338][6],loc[338][7],loc[338][8],loc[338][9],loc[338][10]};end
            339:begin W21 = {loc[339][1],loc[339][2],loc[339][3],loc[339][4],loc[339][5],loc[339][6],loc[339][7],loc[339][8],loc[339][9],loc[339][10]};end
            340:begin W21 = {loc[340][1],loc[340][2],loc[340][3],loc[340][4],loc[340][5],loc[340][6],loc[340][7],loc[340][8],loc[340][9],loc[340][10]};end
            341:begin W21 = {loc[341][1],loc[341][2],loc[341][3],loc[341][4],loc[341][5],loc[341][6],loc[341][7],loc[341][8],loc[341][9],loc[341][10]};end
            342:begin W21 = {loc[342][1],loc[342][2],loc[342][3],loc[342][4],loc[342][5],loc[342][6],loc[342][7],loc[342][8],loc[342][9],loc[342][10]};end
            343:begin W21 = {loc[343][1],loc[343][2],loc[343][3],loc[343][4],loc[343][5],loc[343][6],loc[343][7],loc[343][8],loc[343][9],loc[343][10]};end
            344:begin W21 = {loc[344][1],loc[344][2],loc[344][3],loc[344][4],loc[344][5],loc[344][6],loc[344][7],loc[344][8],loc[344][9],loc[344][10]};end
            345:begin W21 = {loc[345][1],loc[345][2],loc[345][3],loc[345][4],loc[345][5],loc[345][6],loc[345][7],loc[345][8],loc[345][9],loc[345][10]};end
            346:begin W21 = {loc[346][1],loc[346][2],loc[346][3],loc[346][4],loc[346][5],loc[346][6],loc[346][7],loc[346][8],loc[346][9],loc[346][10]};end
            347:begin W21 = {loc[347][1],loc[347][2],loc[347][3],loc[347][4],loc[347][5],loc[347][6],loc[347][7],loc[347][8],loc[347][9],loc[347][10]};end
            348:begin W21 = {loc[348][1],loc[348][2],loc[348][3],loc[348][4],loc[348][5],loc[348][6],loc[348][7],loc[348][8],loc[348][9],loc[348][10]};end
            349:begin W21 = {loc[349][1],loc[349][2],loc[349][3],loc[349][4],loc[349][5],loc[349][6],loc[349][7],loc[349][8],loc[349][9],loc[349][10]};end
            350:begin W21 = {loc[350][1],loc[350][2],loc[350][3],loc[350][4],loc[350][5],loc[350][6],loc[350][7],loc[350][8],loc[350][9],loc[350][10]};end
            351:begin W21 = {loc[351][1],loc[351][2],loc[351][3],loc[351][4],loc[351][5],loc[351][6],loc[351][7],loc[351][8],loc[351][9],loc[351][10]};end
            352:begin W21 = {loc[352][1],loc[352][2],loc[352][3],loc[352][4],loc[352][5],loc[352][6],loc[352][7],loc[352][8],loc[352][9],loc[352][10]};end
            353:begin W21 = {loc[353][1],loc[353][2],loc[353][3],loc[353][4],loc[353][5],loc[353][6],loc[353][7],loc[353][8],loc[353][9],loc[353][10]};end
            354:begin W21 = {loc[354][1],loc[354][2],loc[354][3],loc[354][4],loc[354][5],loc[354][6],loc[354][7],loc[354][8],loc[354][9],loc[354][10]};end
            355:begin W21 = {loc[355][1],loc[355][2],loc[355][3],loc[355][4],loc[355][5],loc[355][6],loc[355][7],loc[355][8],loc[355][9],loc[355][10]};end
            356:begin W21 = {loc[356][1],loc[356][2],loc[356][3],loc[356][4],loc[356][5],loc[356][6],loc[356][7],loc[356][8],loc[356][9],loc[356][10]};end
            357:begin W21 = {loc[357][1],loc[357][2],loc[357][3],loc[357][4],loc[357][5],loc[357][6],loc[357][7],loc[357][8],loc[357][9],loc[357][10]};end
            358:begin W21 = {loc[358][1],loc[358][2],loc[358][3],loc[358][4],loc[358][5],loc[358][6],loc[358][7],loc[358][8],loc[358][9],loc[358][10]};end
            359:begin W21 = {loc[359][1],loc[359][2],loc[359][3],loc[359][4],loc[359][5],loc[359][6],loc[359][7],loc[359][8],loc[359][9],loc[359][10]};end
            360:begin W21 = {loc[360][1],loc[360][2],loc[360][3],loc[360][4],loc[360][5],loc[360][6],loc[360][7],loc[360][8],loc[360][9],loc[360][10]};end
            361:begin W21 = {loc[361][1],loc[361][2],loc[361][3],loc[361][4],loc[361][5],loc[361][6],loc[361][7],loc[361][8],loc[361][9],loc[361][10]};end
            362:begin W21 = {loc[362][1],loc[362][2],loc[362][3],loc[362][4],loc[362][5],loc[362][6],loc[362][7],loc[362][8],loc[362][9],loc[362][10]};end
            363:begin W21 = {loc[363][1],loc[363][2],loc[363][3],loc[363][4],loc[363][5],loc[363][6],loc[363][7],loc[363][8],loc[363][9],loc[363][10]};end
            364:begin W21 = {loc[364][1],loc[364][2],loc[364][3],loc[364][4],loc[364][5],loc[364][6],loc[364][7],loc[364][8],loc[364][9],loc[364][10]};end
            365:begin W21 = {loc[365][1],loc[365][2],loc[365][3],loc[365][4],loc[365][5],loc[365][6],loc[365][7],loc[365][8],loc[365][9],loc[365][10]};end
            366:begin W21 = {loc[366][1],loc[366][2],loc[366][3],loc[366][4],loc[366][5],loc[366][6],loc[366][7],loc[366][8],loc[366][9],loc[366][10]};end
            367:begin W21 = {loc[367][1],loc[367][2],loc[367][3],loc[367][4],loc[367][5],loc[367][6],loc[367][7],loc[367][8],loc[367][9],loc[367][10]};end
            368:begin W21 = {loc[368][1],loc[368][2],loc[368][3],loc[368][4],loc[368][5],loc[368][6],loc[368][7],loc[368][8],loc[368][9],loc[368][10]};end
            369:begin W21 = {loc[369][1],loc[369][2],loc[369][3],loc[369][4],loc[369][5],loc[369][6],loc[369][7],loc[369][8],loc[369][9],loc[369][10]};end
            370:begin W21 = {loc[370][1],loc[370][2],loc[370][3],loc[370][4],loc[370][5],loc[370][6],loc[370][7],loc[370][8],loc[370][9],loc[370][10]};end
            371:begin W21 = {loc[371][1],loc[371][2],loc[371][3],loc[371][4],loc[371][5],loc[371][6],loc[371][7],loc[371][8],loc[371][9],loc[371][10]};end
            372:begin W21 = {loc[372][1],loc[372][2],loc[372][3],loc[372][4],loc[372][5],loc[372][6],loc[372][7],loc[372][8],loc[372][9],loc[372][10]};end
            373:begin W21 = {loc[373][1],loc[373][2],loc[373][3],loc[373][4],loc[373][5],loc[373][6],loc[373][7],loc[373][8],loc[373][9],loc[373][10]};end
            374:begin W21 = {loc[374][1],loc[374][2],loc[374][3],loc[374][4],loc[374][5],loc[374][6],loc[374][7],loc[374][8],loc[374][9],loc[374][10]};end
            375:begin W21 = {loc[375][1],loc[375][2],loc[375][3],loc[375][4],loc[375][5],loc[375][6],loc[375][7],loc[375][8],loc[375][9],loc[375][10]};end
            376:begin W21 = {loc[376][1],loc[376][2],loc[376][3],loc[376][4],loc[376][5],loc[376][6],loc[376][7],loc[376][8],loc[376][9],loc[376][10]};end
            377:begin W21 = {loc[377][1],loc[377][2],loc[377][3],loc[377][4],loc[377][5],loc[377][6],loc[377][7],loc[377][8],loc[377][9],loc[377][10]};end
            378:begin W21 = {loc[378][1],loc[378][2],loc[378][3],loc[378][4],loc[378][5],loc[378][6],loc[378][7],loc[378][8],loc[378][9],loc[378][10]};end
            379:begin W21 = {loc[379][1],loc[379][2],loc[379][3],loc[379][4],loc[379][5],loc[379][6],loc[379][7],loc[379][8],loc[379][9],loc[379][10]};end
            380:begin W21 = {loc[380][1],loc[380][2],loc[380][3],loc[380][4],loc[380][5],loc[380][6],loc[380][7],loc[380][8],loc[380][9],loc[380][10]};end
            381:begin W21 = {loc[381][1],loc[381][2],loc[381][3],loc[381][4],loc[381][5],loc[381][6],loc[381][7],loc[381][8],loc[381][9],loc[381][10]};end
            382:begin W21 = {loc[382][1],loc[382][2],loc[382][3],loc[382][4],loc[382][5],loc[382][6],loc[382][7],loc[382][8],loc[382][9],loc[382][10]};end
            383:begin W21 = {loc[383][1],loc[383][2],loc[383][3],loc[383][4],loc[383][5],loc[383][6],loc[383][7],loc[383][8],loc[383][9],loc[383][10]};end
            384:begin W21 = {loc[384][1],loc[384][2],loc[384][3],loc[384][4],loc[384][5],loc[384][6],loc[384][7],loc[384][8],loc[384][9],loc[384][10]};end
            385:begin W21 = {loc[385][1],loc[385][2],loc[385][3],loc[385][4],loc[385][5],loc[385][6],loc[385][7],loc[385][8],loc[385][9],loc[385][10]};end
            386:begin W21 = {loc[386][1],loc[386][2],loc[386][3],loc[386][4],loc[386][5],loc[386][6],loc[386][7],loc[386][8],loc[386][9],loc[386][10]};end
            387:begin W21 = {loc[387][1],loc[387][2],loc[387][3],loc[387][4],loc[387][5],loc[387][6],loc[387][7],loc[387][8],loc[387][9],loc[387][10]};end
            388:begin W21 = {loc[388][1],loc[388][2],loc[388][3],loc[388][4],loc[388][5],loc[388][6],loc[388][7],loc[388][8],loc[388][9],loc[388][10]};end
            389:begin W21 = {loc[389][1],loc[389][2],loc[389][3],loc[389][4],loc[389][5],loc[389][6],loc[389][7],loc[389][8],loc[389][9],loc[389][10]};end
            390:begin W21 = {loc[390][1],loc[390][2],loc[390][3],loc[390][4],loc[390][5],loc[390][6],loc[390][7],loc[390][8],loc[390][9],loc[390][10]};end
            391:begin W21 = {loc[391][1],loc[391][2],loc[391][3],loc[391][4],loc[391][5],loc[391][6],loc[391][7],loc[391][8],loc[391][9],loc[391][10]};end
            392:begin W21 = {loc[392][1],loc[392][2],loc[392][3],loc[392][4],loc[392][5],loc[392][6],loc[392][7],loc[392][8],loc[392][9],loc[392][10]};end
            393:begin W21 = {loc[393][1],loc[393][2],loc[393][3],loc[393][4],loc[393][5],loc[393][6],loc[393][7],loc[393][8],loc[393][9],loc[393][10]};end
            394:begin W21 = {loc[394][1],loc[394][2],loc[394][3],loc[394][4],loc[394][5],loc[394][6],loc[394][7],loc[394][8],loc[394][9],loc[394][10]};end
            395:begin W21 = {loc[395][1],loc[395][2],loc[395][3],loc[395][4],loc[395][5],loc[395][6],loc[395][7],loc[395][8],loc[395][9],loc[395][10]};end
            396:begin W21 = {loc[396][1],loc[396][2],loc[396][3],loc[396][4],loc[396][5],loc[396][6],loc[396][7],loc[396][8],loc[396][9],loc[396][10]};end
            397:begin W21 = {loc[397][1],loc[397][2],loc[397][3],loc[397][4],loc[397][5],loc[397][6],loc[397][7],loc[397][8],loc[397][9],loc[397][10]};end
            398:begin W21 = {loc[398][1],loc[398][2],loc[398][3],loc[398][4],loc[398][5],loc[398][6],loc[398][7],loc[398][8],loc[398][9],loc[398][10]};end
            399:begin W21 = {loc[399][1],loc[399][2],loc[399][3],loc[399][4],loc[399][5],loc[399][6],loc[399][7],loc[399][8],loc[399][9],loc[399][10]};end
            400:begin W21 = {loc[400][1],loc[400][2],loc[400][3],loc[400][4],loc[400][5],loc[400][6],loc[400][7],loc[400][8],loc[400][9],loc[400][10]};end
            401:begin W21 = {loc[401][1],loc[401][2],loc[401][3],loc[401][4],loc[401][5],loc[401][6],loc[401][7],loc[401][8],loc[401][9],loc[401][10]};end
            402:begin W21 = {loc[402][1],loc[402][2],loc[402][3],loc[402][4],loc[402][5],loc[402][6],loc[402][7],loc[402][8],loc[402][9],loc[402][10]};end
            403:begin W21 = {loc[403][1],loc[403][2],loc[403][3],loc[403][4],loc[403][5],loc[403][6],loc[403][7],loc[403][8],loc[403][9],loc[403][10]};end
            404:begin W21 = {loc[404][1],loc[404][2],loc[404][3],loc[404][4],loc[404][5],loc[404][6],loc[404][7],loc[404][8],loc[404][9],loc[404][10]};end
            405:begin W21 = {loc[405][1],loc[405][2],loc[405][3],loc[405][4],loc[405][5],loc[405][6],loc[405][7],loc[405][8],loc[405][9],loc[405][10]};end
            406:begin W21 = {loc[406][1],loc[406][2],loc[406][3],loc[406][4],loc[406][5],loc[406][6],loc[406][7],loc[406][8],loc[406][9],loc[406][10]};end
            407:begin W21 = {loc[407][1],loc[407][2],loc[407][3],loc[407][4],loc[407][5],loc[407][6],loc[407][7],loc[407][8],loc[407][9],loc[407][10]};end
            408:begin W21 = {loc[408][1],loc[408][2],loc[408][3],loc[408][4],loc[408][5],loc[408][6],loc[408][7],loc[408][8],loc[408][9],loc[408][10]};end
            409:begin W21 = {loc[409][1],loc[409][2],loc[409][3],loc[409][4],loc[409][5],loc[409][6],loc[409][7],loc[409][8],loc[409][9],loc[409][10]};end
            410:begin W21 = {loc[410][1],loc[410][2],loc[410][3],loc[410][4],loc[410][5],loc[410][6],loc[410][7],loc[410][8],loc[410][9],loc[410][10]};end
            411:begin W21 = {loc[411][1],loc[411][2],loc[411][3],loc[411][4],loc[411][5],loc[411][6],loc[411][7],loc[411][8],loc[411][9],loc[411][10]};end
            412:begin W21 = {loc[412][1],loc[412][2],loc[412][3],loc[412][4],loc[412][5],loc[412][6],loc[412][7],loc[412][8],loc[412][9],loc[412][10]};end
            413:begin W21 = {loc[413][1],loc[413][2],loc[413][3],loc[413][4],loc[413][5],loc[413][6],loc[413][7],loc[413][8],loc[413][9],loc[413][10]};end
            414:begin W21 = {loc[414][1],loc[414][2],loc[414][3],loc[414][4],loc[414][5],loc[414][6],loc[414][7],loc[414][8],loc[414][9],loc[414][10]};end
            415:begin W21 = {loc[415][1],loc[415][2],loc[415][3],loc[415][4],loc[415][5],loc[415][6],loc[415][7],loc[415][8],loc[415][9],loc[415][10]};end
            416:begin W21 = {loc[416][1],loc[416][2],loc[416][3],loc[416][4],loc[416][5],loc[416][6],loc[416][7],loc[416][8],loc[416][9],loc[416][10]};end
            417:begin W21 = {loc[417][1],loc[417][2],loc[417][3],loc[417][4],loc[417][5],loc[417][6],loc[417][7],loc[417][8],loc[417][9],loc[417][10]};end
            418:begin W21 = {loc[418][1],loc[418][2],loc[418][3],loc[418][4],loc[418][5],loc[418][6],loc[418][7],loc[418][8],loc[418][9],loc[418][10]};end
            419:begin W21 = {loc[419][1],loc[419][2],loc[419][3],loc[419][4],loc[419][5],loc[419][6],loc[419][7],loc[419][8],loc[419][9],loc[419][10]};end
            420:begin W21 = {loc[420][1],loc[420][2],loc[420][3],loc[420][4],loc[420][5],loc[420][6],loc[420][7],loc[420][8],loc[420][9],loc[420][10]};end
            default:begin W21 = {loc[1][1],loc[1][2],loc[1][3],loc[1][4],loc[1][5],loc[1][6],loc[1][7],loc[1][8],loc[1][9],loc[1][10]}; end
        endcase
    end
    always @(posedge clk)
        d<=W21; 
endmodule
